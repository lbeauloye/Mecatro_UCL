    Mac OS X            	   2   �     +                                      ATTR      +   �   o                  �   S  com.dropbox.attributes          com.dropbox.attrs    x��VJ)�/Hʯ�O��I�L���ON�Q�R�V�ML����%����RK��2��B��(�$���b�� �LsC�r[[���Z �(2

�!�WJ>�     ��ˡ�