    Mac OS X            	   2   �     +                                      ATTR      +   �   o                  �   S  com.dropbox.attributes          com.dropbox.attrs    x��VJ)�/Hʯ�O��I�L���ON�Q�R�V�ML����%����RK��J�
o#K#7�P�tw�<�,��@[[���Z ��

�!�WJ>�     Ѭ��ݟ