    Mac OS X            	   2   �     +                                      ATTR      +   �   o                  �   S  com.dropbox.attributes          com.dropbox.attrs    x��VJ)�/Hʯ�O��I�L���ON�Q�R�V�ML����%����RK����2�Ϩ2�R��J�RW}Ggӈt[[���Z �Zb

�!�WJ>�     ѻ����