    Mac OS X            	   2   �     +                                      ATTR      +   �   o                  �   S  com.dropbox.attributes          com.dropbox.attrs    x��VJ)�/Hʯ�O��I�L���ON�Q�R�V�ML����%����RK�%��㢈�DK#7�0ϠR�SG[[���Z �?9

�!�WJ>�     �8��Ċ