    Mac OS X            	   2  U     �                                      ATTR      �   �   �                  �   <  com.apple.quarantine      S  com.dropbox.attributes     k     com.dropbox.attrs    q/0083;5c851a5a;Safari;84C2A4D2-7C4C-4732-A127-443F1530B6AA x��VJ)�/Hʯ�O��I�L���ON�Q�R�V�ML����%����RK�%_�$� ��t�tG��� ϴR�мt[[���Z �?�

�!�WJ>�     �����