    Mac OS X            	   2   �     +                                      ATTR      +   �   o                  �   S  com.dropbox.attributes          com.dropbox.attrs    x��VJ)�/Hʯ�O��I�L���ON�Q�R�V�ML����%����RK�%�3�Ĩ��$W�
�J�r#��r[[���Z ��$

�!�WJ>�     �n�ځ�