    Mac OS X            	   2   �     +                                      ATTR      +   �   o                  �   S  com.dropbox.attributes          com.dropbox.attrs    x��VJ)�/Hʯ�O��I�L���ON�Q�R�V�ML����%����RK�%�
��Boc�Ĉ�4}}�@�˔r[[���Z �7�

�!�WJ>�      �ݍȽ