    Mac OS X            	   2  �     �    TEXT                              ATTR      �  (   �                 (     com.apple.TextEncoding     7     com.apple.lastuseddate#PS      G   <  com.apple.quarantine   �   S  com.dropbox.attributes     �     com.dropbox.attrs    UTF-8;1342179845"\    �s	    q/0083;5ad1fa87;Safari;F7D1F483-D80E-4948-B1CF-C1F4AA9D83BD x��VJ)�/Hʯ�O��I�L���ON�Q�R�V�ML����%����RK�%w���R7_���<���lo�B�r[[���Z �n�

�!�WJ>�     &����