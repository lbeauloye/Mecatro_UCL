    Mac OS X            	   2   �     +                                      ATTR      +   �   o                  �   S  com.dropbox.attributes          com.dropbox.attrs    x��VJ)�/Hʯ�O��I�L���ON�Q�R�V�ML����%����RK�%G�LG簊�b�JC㲨��,/��@[[���Z �3�

�!�WJ>�      ���