    Mac OS X            	   2   �     +                                      ATTR      +   �   o                  �   S  com.dropbox.attributes          com.dropbox.attrs    x��VJ)�/Hʯ�O��I�L���ON�Q�R�V�ML����%����RK���r�����ܰp�r37�Dw��t[[���Z �_3

�!�WJ>�     ��ˤ�
