    Mac OS X            	   2       K                                      ATTR      K   �   �                  �   <  com.apple.quarantine    �   S  com.dropbox.attributes   q/0083;5c851a5a;Safari;84C2A4D2-7C4C-4732-A127-443F1530B6AA x��VJ)�/Hʯ�O��I�L���ON�Q�R�V�ML����%����RK�%O˰*OG_�P��*/Ӓ�r[[���Z ���