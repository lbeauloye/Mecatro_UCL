    Mac OS X            	   2   �     *                                      ATTR      *   �   n                  �   S  com.dropbox.attributes          com.dropbox.attrs    x��VJ)�/Hʯ�O��I�L���ON�Q�R�V�ML����%����RK���� c��|�|c'���bS�@[[���Z ��	

�!�WJ>�     ����h