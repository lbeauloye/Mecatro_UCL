    Mac OS X            	   2   �      �                                      ATTR       �   �   S                  �   S  com.dropbox.attributes   x��VJ)�/Hʯ�O��I�L���ON�Q�R�V�ML����%����RK���4#�`��0��(�������@[[���Z ��Q