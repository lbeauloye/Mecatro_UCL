    Mac OS X            	   2   �     +                                      ATTR      +   �   o                  �   S  com.dropbox.attributes          com.dropbox.attrs    x��VJ)�/Hʯ�O��I�L���ON�Q�R�V�ML����%����RK��t?�PǴp�r#7���L�4Ӭ�|G[[���Z ó_

�!�WJ>�      	ӟ��