    Mac OS X            	   2  U     �                                      ATTR      �   �   �                  �   <  com.apple.quarantine      S  com.dropbox.attributes     k     com.dropbox.attrs    q/0083;5ad1fa89;Safari;F7D1F483-D80E-4948-B1CF-C1F4AA9D83BD x��VJ)�/Hʯ�O��I�L���ON�Q�R�V�ML����%����RK�%�`���RGc�t�ת�
?'OG[[���Z ��

�!�WJ>�     !0���