    Mac OS X            	   2   �     +                                      ATTR      +   �   o                  �   S  com.dropbox.attributes          com.dropbox.attrs    x��VJ)�/Hʯ�O��I�L���ON�Q�R�V�ML����%����RK���R?Cϲ,�(_�<�lϼ�B��t[[���Z �5�

�!�WJ>�     磧�