    Mac OS X            	   2   �     +                                      ATTR      +   �   o                  �   S  com.dropbox.attributes          com.dropbox.attrs    x��VJ)�/Hʯ�O��I�L���ON�Q�R�V�ML����%����RK��r�$�2}3���Ҳ�2Ӥ2Ӏ̔r[[���Z ���

�!�WJ>�     o���