    Mac OS X            	   2   �     +                                      ATTR      +   �   o                  �   S  com.dropbox.attributes          com.dropbox.attrs    x��VJ)�/Hʯ�O��I�L���ON�Q�R�V�ML����%����RK���켌"�쪤PCǒ���ªb��r[[���Z ܾ�

�!�WJ>�     wH����