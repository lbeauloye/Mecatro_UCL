��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���QΠ�F�p��������m܇�+�˺7�)H!A)=8N���`'��N���K"��}�m�X��J� �e}�<���]���*`�F�Y�EF�9�j�ChT�1_ ��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �&����y���^ �Aq�&�����Ղ8�~��kD3~�bVwv'4�,�\w3-�P�^1G��8jH��|�Sq���� ��`�h�r�%1\��Tjk��qJ�T�"��]ۓ��P�Ҫ{�����`�w��c Mq�`CΦ<'c�>�"bxw]�؝ϳl�Yya�e�=���cq��oc~���25�ԭ���I����Dj��b`�V=�}�\�ڸ�E�y  ���N#w�������!������v���Yb>3������ō�c�Ҵ�	��C���g�y�B�W��0�WB=Ai���[Q�Y�q�.l��zDl�y���(�Ē"$��m�?-�i=�D�D&,>z�{g���觪sp�c�`X[�K�֤�M�]��ٲ�o���\ 	���Y�_�;J�LN!�Im@_�/oo�¨�m���O$w'�'i]��:0��9��^��b61�_N�!�f��-���4�f^���EI'`�[�nod�/�^��0�<��TT�����C��ɀ2x<kk��c�e�Y�@*�k�m�ݕ��w��C����}�^_��4"k���d�|��� ]�E��v>O�GP��	�:�a�v@X���{��.KTU2=�蓠�~0�w�"��e�V�y�;���lQ|�8�v�h�v�� �oh�ē���آ>���n+�o��IѪ	w����g���tTu�@���gtT�)�J�V�^_D���8�T}��ve�rT@�>�v�ϵ��K�{>ǎ'�GYބ���y~8�pn����P�����(�Os*��>1�㤪e8�+�1F�E�d��q*�Mp�x��h�6��H�Bs+�t�4<<�sn��<���¼a:��NB�ϣ	?F�	��|?��'5a��S󌼟�W��p?X!�kP�&ݱBġ�U��9v$��e�)�M �?��wh`+��b)�f%�ժ���Ǔi���m�+�J'�{�W��9��π�`��|&1($�cӢ�-��Ω5Z�Jɗ
սB��1-\��#6?ޅ\f�q>�pu�,qK�a�4���O"s��[L-��84��_RigٜML}�:9L�.�e�y�7E���C���F�9�]9�O�fG����cu��0$���j2�}��P1�%~aW�h�`�Z��cL�;��}����c�[����9�
�%��F��y B�]�Rkf�S���(?:�y�����B���R��C^-�b8^��٤�4��՝kC�����{e>]�	��X����Ue�;/P�"�1�]�����/Vp�&MqH8�F��O�cLb�?���?��f2^���4��7�#� 8���Q��JGG=����o�z7#ڵ�Lݨ���~8��:��kk�)�XC���.�"8H�R,0����_�R�F��#��=F��)�Ab�#�Sq=�*u��Ša��M��p��8>B�g�h��I�R���*Fg[qǝU��I���Xu���g~9�z�a��/Q!���_���"P���ao�b�A&�<q����Y{u�a��
�������[�_������
��ӟ�G����Q�f~�,�&�;7D���bL��ٲhF�L��cf9އ�(�.v�n�q���\*������'��ɦ̨�N�n�2Z}�`��e6�v�Q����O������]�Sӵb�9o���z�Q���7a�Lr�]�Wst��ę-lqć��c�&tP)�⏎C�c0��"
g�Z�T�\��I+Tn<�*�liE�ҭ�&㡆:C�+yբ��7e��I��A�tɿI�5�־�c�ޮ�e�&�i.��d@����秣��� Db�Z"l��_?�[����}�]�v�a��~��?B�&��å����\d������'�V=�@d)?���� 1�+� �Щ�dY2p8��"��2t��iŊ���t����R��ZutFf:�j�J҇��0��Y�t~N�5�7>;�0�.a��J��G���䴘D��]����P/_���9G�>�&�oJp�Ӕ�Y%����p܄Ǚ��	�A*�	=�I�[��c����a�Ӭ�b��s:��P:���0�P���1~Ŝ]+�ājKb�yNw��E��o�u��W��N܃���w%M���ߓ�z1)D�I�2�j&&H�j2�����Q&)#�@!h��0�|S�0,�g�b����1�0H�4����)WC���"�Z2k_�U�6<thN��[.�*����֒ʔ����w�)��,��\���c�;Yi�l:�9F����bl��F�Ӂ��	o�����R�]q5\������k?]�BC&*y�97Y��o�b0J<a����;�eq����8�0���	�ZyS��;Z��� �2��_�ƌ�4���[QZr؜}9o�	�ʥ�ˁ;$?���m���p�t���>	���Q۪|ǳ���в���Uط[{8�E�Nw(tM�����`�`W�d��``�E7	[��u���K �|����2�T���^e�������gE[���	�n��GU���~�a�L54���;�-	Ii�o��f�＂�Cv���v�y�K���I�w+��¾[3K�҂:/��$m�b0��b@YNE�l@�M��/fyZKJ{Z!����)f�f�"��O#��j4�w�I8���gg� D����QU�������
|.2���j�4����-ۡ�ν�� ��-ۜ"-�ͳ-�����7FJri�(�g�+����9�;�^�b�D�v���X���
��Es��<3�%�Z��m:W�H��|=d�p�$���?/+�,���c��Y���0)q�n�#MJ���Zu�>��t��YI���O2����2Tu����L�
y� �WFZ��$��U�&��(���sK_MO���q�^V���D������s,�.� �L��]B~����4!	θ;RV��d!8�#֭8ʮ-Q{P~�"�?%�VU%����cmPѯ�JF^a�W���vM�?�!�gv�Yt��7����"�=�.����NwB{�	�V�U���(�TP��Q���ٻ�� ʔ(L�]�"e�V�~e�z&&C,0g�=�H���*���&#�3U���k��	���R�8>)��/���9B��\N��ɷ�~�f��}ⳘPB��:�0_������J����,��6R`���j�,M�E���bЉg̟$v��D�c#��W��mk�Q�t�����>!GQQ����Z�H!#�:�f$�/������hE�AW?6'�5�˽K��~t��7y�/�4�#�x˸2���$4�����aHN4����yWv[Ƅ�א)E����ۣ(~[���"��ϒ1�3έAI�����#ݚ{\j�j_��J>QɹoC@�����}��/sY**mη��׸�+�y"o"v�o���W�Zf�͝�'�c}-*�|0�n�ō !k��J�";ƹ�h�������b��g�����1[o�<���~
+�oP�*���ѧ<��i���dA�(PY��]�U��h �|>N���:[k���!���m�B!f@��Z�C��4:?Ҕ+��� �ݿ��x�B͕� �֧^��U���pp;�,�!��-̷5Z5�	�m!'l�7Bf��d^��uu�kр_V2��>� �N��]9�!��E@6�a��)ǸFi~�k��NpsRH0f��戹>r����;�=�Ĥ���;9�S֚��1�W�7��Ch6�$���1b��w����D��N_��O00��W@Z�\n����(S��^��F�r��7ar.pp��~#�o��0����g	�:�IS �7��e^+N�@��.�w{f�C6)zP���R��Á,c�-�N�}�u�\YD��C�-�|�42��G�]x��vc���̴��ڦ�7��FK�
���En�� 맶 ��X�J�ǀ��hda*�M�l���Pwr
\P�}���|kQᅻ���*E��n��R�3he����������is\�'I�܉hP*Y�Z�M�I&�K������;�Sv��+�9l�~#���.���%՞ק�s�M��['e6<��C�+p0·���A����?�(�2;��F׽��tR�\޲^������E�N����.��u��*�`gӺ�@���#��N� g��6Ƿ�W�g�d����_���(%�G�ȿ�K�BU,.1V �R��xي���~�x5׼����/B��p\o����k�}�O�3�C��1�P���{YA��%���X@�HF�{vV�F&�/��Jfk�u�F�w���a�A*�W��JE�g�qN2[�:���I�+�����@�Tj�.Jl !�c-x Tdt�B������9�V�(,T��IܧP������JJA���
5Ye����hVH��m�d�����a�v��	�����Zt�Pg�U�C|N���S�؏��3�M���F?7�]fT��;@�Z���`����$��n���?SmY(G��v���7���G��u)��.u�ܯ�`�����l- 6z^�_�ZLW,�Ĥ'��Q��h�p--�@��uS�Z�:=]�BFs�ډ-g (���T�z m���눒e3��4,\��'"�foG���N~�|�@�uG�CZ���vh�-]>�Zi|�4�]BsZ���與HGH�8�:&��1A��c�fpPԬ�ʯ?�$vAD\�Y��b��N
?Liʿ�<:��/H�s~|�X7�B���YP��,l�����kP6�+�)��y�g������w�>R�F�Qꀵ* H���
����@Б���w.1��e�Cwѱ+1U)���Ǘ�Ε���`СWt*8|��f��zԦnݢ����fK9�&�{>���)�����Ꭷ��M��p���a� �زla��S9W�j� !q(��~����SR�ϔ�B����|�h�ПRk}Ϩ�؛�0K t�(י�E�ܰ�fӓ���g�K
��-jeU�����/�2��׮J���%���9��wB^xO�左�UM�ʶ��Q����$$����ʠ��ٵ��3xv
ϳbCW�Xu�2w�#�.=®pP7[���±�J���l��ܺ�����d�-��r�I#:l1:��]�X;��:H_�Y�k�'��(z��`=f�Y(��KT��v����y�{���0�������Hp�c	h���O�Z�2&F�żG:l��J�h\o�q1P<�"�}���9��-z��,D���@��R�k|0Ϧ�ˢa�Y)Sc�|p���1���#f譜��kc����z�Ώ���-��[�|u�a���%��|�	Eا'�9!ݐKtS��F� ar�&�.����}�9�f������������]�M��r��[�%$�C�X�<=ғx	}Q��q�<#�z(}��N�!�z�2z�u�
�x���UQR���N��Py�d�U�v`��%g�;G�YgNa`WK�Yo��$ЌqCTi~F�5���DU9J���(�w&���ݑwݙ%�O\����v�-5$1���H��U���i�Fk���:��q)�\q��5)��V|������2 ��}�ݥ��(�K�bH�1�h�ec�odE���p�
�Ȩ�u�s��`��z�##�U�?�nZ�؍*F��0it޹\iPi�j� TD4�"�����p9q��5�ᠪ�q"b�~�D�y�1��_�|$ ��SN�Ew|���:��a�9�½��m�p�!�=^��u�4uk�E����7$�P�C�ކW��U��$�oG����t�:�HW{\��D��1䱢Ǣ����}W�}�R���N�3��Ixgć�jDcC	~V@��%k�9o7���-rm�x%�]p�O�]�;Q2O`0�0C5hl��v���o.|~̝z슈��٤�I����X���YiN���C��kse���p
��-�q2��8b$�1�lCKNߴ���'�*��}>�k����]z��OE9`u���ۻBFw��z^��4҇g�sZ)A��ťϢg��7�9"h�x��u`ܾI�z�������=�*��i����������2ށG^/������s�4b�p1{��C�:�*�H�U��H�v��<�E�|0lc��t2��>�L*O��ݹ�%%��V�j�G�}9�*S� ,RbK�"F�o~l���2j�]���s�؃��]�7��>#�+�� ��P�Z�s�����80r��	��C�o��<�����v�0�?Ѐs<�wrJKa�l��#�%H�W�x����*�:��f��Z�GN�&�ՌY�M%��e�����b�:��p�[c��B/��C�@�Hޮ9�}���R@���[��ƌ�ry��L���"��im�B��*	A�����U�bl�^7B��K�W�0yb@����2�3�Y�K2,�K9b�8�>��J �t�n�X�l�X���E�VN�d�����g!B���Rs�I����'�I�k�5��̔��lk�bPoj5ɟV��e&�~V߲G��U&u�����0��Ğ
�.J�r:�;j;G��	�wa�TJ�f����2����[�/���'�����uCdg��4J;�ͨ��{�<L>ƍ��\'DH�Q�[14KJl��`���Kcl�	 ŏ�:J�����g4���h��x|�j�f��N+��a��W͌ M�+��
K:cX��H�(ujq�O��(�j�N�����ّk�mA����D$��[�2m<����a-WMJ���lٕeZ��	Bm�1k<�����nx|�ɯ
��Z|*��7�n��8��$F��
/.^�:2PM�E2zU݀Y��4:�YapoD��Ĝ�7������| g�L��%���D�Վ����ઐW/ly��ꜚq�{NB���jY�A��*�4e�!��_�Go��F����DC���UF��0�@ 7�S����ȥ(�4uI��G�v9�������V��auA��c� �mc@��|ԑ����w�<ݷ�L�eI��7��9�s���S�FU�PZU�0�=\����Z�+��P�q�J��x��,�T)ڲ��q;�~����۵���=
���)y~�!�S<?����u���F�qP7T��I$�I�J�g5~�3\v&����)�$Ÿ�@ ]�O�$~<۳ �`@6 ��D^ɣ���E$��*^8Z��ڽx%pi���=F����gp���*�Y�*@LN-���� ���EZ��b̀�;���G��� ©m[m�������x?Ĩ��󼈕�dhm�e�F�ĆsT�!=,����e�;̅��o��6��'xk
�}%��z�럓�^���S�,�	�O<��k�BL	ʀ��P/,sҏNL�����&C��+����������z��v�N��������V��Nt�����pTP,��3�{�|+H��86��(K��r���˻���
3,�8BeKi���8c�՟8�A��X������_]˔ X��x��s[8�x���
0P&�z��A|����*�i�7�W�pW^2��s`���e�� ��E����Yjb�[,ز
���i_T����Ht9�,�3/1K��V�j1�No?���(
��f���ɭ����%�\�k�n���ϊuU���w'��O4�5Xm=a�A�ؤ��B?����u��^F�me�z�ŌJ�G0���������ʃ���V^?k9j
��f��0��S]�S�y8�=�z�(}���␐�{.��PK�%6��9m٬x����xk��)�!�j���R�қM=�0�+��=b��G�֫'u*�<\.pI��)ͦ����uŧ��~��/tj�'�P�Ht��C�lM C=�PFa�S���Ⱥl��-?D=!���]����:��� 6�hIѳ��ȁs�{���/�A�P睢N�Tgk��b]
���%���Xu_��}K��0'*F%�!~��a|�+6_ }��u��Cy�"�[<��r��a���FON�����g�u���ǆ��e�?8�vF��=ErA��T�z���F��rfڑ,�ڣ`���:H��{��kr�L>�v9*'<�T�)7妍i��m`+��K���*:�!��7A)�[�OVu�<w,S�O�8�Z�ꠝ��ǟ�zK�)5b�6(oJ�֭������	>ݰ��UG����3��u�85��2%�ƌ�,�0����z�:�l�(�-H�>a0&q���a�
��附���c[K<��F����v��؝��{Q>q�S�@Km���7T
)0
՚7��I�E<�-�]�ʩބ��L�Y���O�ְJ"��	0�QZ�%1�:�Z�7��k�j��p�f
���Q�F}FI|6�"fg^�����
�(���oI�T�E��"�7tPV��@�0�=*���x��[:(�oObl�H�#sN�9(II�!��a|�X�5C�-�o���}����G�ɧJ��G6���/���6�{M�{Jb�����*'��9KU��e�-�ۭL���>l)�f�Cd2�3i"H��u�P��������u���z�F�l]��T��ؠ^��G��B���W�@0�����cN�͋��fp�f{\�#%��E��*�)u$G�Ɂ�e�i�4Kڰ.&�y���w�mşђGV�=����#��#W�I&��O���}�	d��iv6<?6�8��8�ެ�s���!x��9#=�c�Ϫ47����f��%�7wi���BAx�k����x�$�`�pt��ř�0�o�R�]�;06[�Uꍑ B��h爡Xv{9mqίr�����I�_FJ��L���$���ki�#c� ��0<N�r��N���عE�6�����I	�<:�y.v&@�#�2�X���:��
��"�ֹ
z��m* )��:�)�;����\�GxvP�yl?��r�=�%l��ɪ�w��5jt|� c����턃{,%�+v<�����6�I�s�u��W'n�2�&��ߞ����R9y������*o��+��&��6�];_lB��(�X��.!F3�8�vy�;g֑�[����3�t_I!�u��+�Q,90������V"O"�hei���٭Aw����naH ��O�7<CPC
H'ں�<4�� Ӳ�Qy����|�E/�&\��G��
�|��Ҕ1�����K#�~�a?���E��i	s��� z�:@��~{猱g���/����&¦*���� �j47�gcv�x��O��!�f-.X�o���Kpf����%~��AҮ�xC�DJˣ�2V���sZ���+�@�40�R�df�w.�wu�ŭ(���2�}ѕ���{�u]�?��@f8�_��z�(j�rJ1����nm���œ9�;�<l���zS�������~��B��a�J�1����|���!Dm�z2 H���XaAV�)�\���f�������R?L��J����3�H,fF�S�Q�g0ӛe�]e9럻�w���<wq].+SW��0�&?P{��;��%	}�)�(��b;M1L�<؊;7�k�S��x�Ǎ��ۺ�_E{�.�� =����j�h�G�M�g��p�P�4��`�%0Ȓ}�	�E�êI�	ѫC��0��):d=��?���V�gOM�	9�cJ6%)C	�����E���%X0g|�m��q�t�;�y�׷Y�(�)��G�池��������	?j��`P7��&B�*@��R��?�i�st����΅�����uȶ;4ĵ)�a?u�X�v�r�kxl�Ig�K��ɺ���D<*?xˇ� Յ�ᮖ�!�0�	�]��Y{�tz�L%������[��xG[t-C�IHQ���.vGa� ���+8�K��o�閁���ǚ��s[��D�pڜ>oDrD�r/���.��80��X��	�O���
��a�)	�~�A5�������B+��O��ieD�߂�|{�5H��h��e��A�q����uz�����UE�9;�0�r%�s�[��ìW��.��!����'�d�l!,��!-������{Ҿ;�yh�/Wx�PXu�}��]��!@� q=W�V�A�( ��9����[����i�>"��|�H.4�;�oҢ�/� ��{4=r@Y���MreX?�S�q���=��I���%1}�R�`�v=�_!
!�s}�@.@��m��D���z�V�q�j���̶���R�+ �]����C���4d�m9w�^'� ~�gk_̅x�Gr���+�FF��z�e��?��?�N*� ��\E7��'?�%���x�v��|ו��!v��}\ *n�+�aV���A������7�<8��ߑ^���u#Ziƛ�q�>(e��S*��0��G�.��q�w��UdL7đ���?����+�Q�Y]����8���&���=ɑ��@��8��Cs;��c_�!�hI�eV
z�:�^�6a8��5,�Wa%��ŵV�4��4n.`�e�xkݻ�EΪp�����M�{J�*R�ɗ�l9��΋����gt?2�]�Y�����	]���gNnc�FE������め�$jF��?�-�Z�.b{�<Mg���hr�Zq�����A��%Az�@�^`C�m�)��E�=s�>�;K�5y�r���=�S�
��J����L�h�<a(���؇��e��jO��\����5��YAk"0�6�=Ie9����������|��A�-]G!8+Uߐ�#v���k+3Y�<�,�i�����MG�)@����s���� ��2�2������Ջ�,Lkc���$ S=͈N�I�����G�����q���`f�ug&R-�P���ׇP3^(�f�HK(�m'A�~*�eA�os$mz�	v�	��,A�b����~�Zge��y�eܥON���X^�e���}ʀ������B�H�t��/bLwQ<j���x��*�/���\�б�� ����l�6�,d���j)�SaS�"�}�E�-�9f��[��6`�E�j"X<�Q���C ����z�:�����Ӣ]�2U�U
�h�sv�����n"o�dó0r�o��aO?�񃐓J���t�~5����!�<��"NT�����'���߫8����Y�~�.�I��o�;^���Z��ƸW�r�z�3�������THh3Q�I��Е$�%��,k9�fd� ��uV�����>H�\B����9"%s�i����o`�Xh��=��,ʔ�4����K���n^��4MJ�phU��Yv)y���W�Y q#��s�Gs-;iP��fz��T!!�=�T�8��|!��i��h�LS��sN�쌧�ӛ�e �7��r{�څj�M���hC�nB�|�^&y^�ۙ�4(A�G#����1��tV0'�.	���V��u(u��ab?eƥ.D�z���d�'�j��3��
D�����:ż��3\�[zW��"z�ٹ�lY�G��/�ݞ��rn�a���w���W&l��?�l(�"�qX��WV�������z�	\�Bt��}��1?���
� �E{A��xy
����]Ct�:�rԬ�VT���K����Fl�����������]�u6� �hvJ��Q'�}���[��Zo��h�Z�[ {=�����&�Y$B*���� �:ጼ�;�n���Y`�e���u+Ŵ��k���p�h�0�m_�叇�@'���4��O���˷�7�WѲ
.:�F�%�.�"{\�e>*�/�mt�$��sÒ�ɹ�e�.��Ӗ���r�΋�4��2���X U�f{*W�2>���c�}q0"��g�c���U�8k�=�ٕ��V"�Ń#}S��}� �>*>Ob��<\����0}85��%D�qA��}^�9��J��5V�����*�M3���=�#ŸB��|����kL�~s.F���<O(���.Ϧ���K���������W���"��:�\ӌzanQ��"h]a�V�� $K����0i�W�I���k���3k�ߟP?������s����&��n�|3r�يD&��6c��V Y����'E��4�vu�1��o&�m?6d��	��ԙO0{�2��_�����H�<�C	�p-���9܁����Ո?�)��h�<Gl�^.,G�ؓǫ"����ىJ} �yc��p��;RiѶVq�����.Y��+�9����ݶr�9�Һ�U�E��4k��?�ϖ94�"
Z,�v�Zf�I%�������HN�9���0����@W�gb�yz���|�#�����1]� ��� ������	rW/�$Z��(�lU�<)�n�
���C�GW (�g�1��L�z��<&��$#�K�H����dV�WJ�H���?j��r(�eU���П�����DR6�($�@����ʁr��LK�1�T��Bi����I'�K��hs�՝%=���J���Q��׆y;�}�T}��)<���rg�Ke��+������&(s�΍9ɬ�dM���^�����E�s��Ӊ[�V� ��`��k�������H��J�ؔ�v�T��:[��%Mv�@.<�m���1��5���R���Q�xj[��R8�dUeظ��_�$���.�ע+��/���Utr�/,W�f+��	CB;�� ��K�ˉC\ɋU4V��Ze��e� ��F$�!-�0�G�����wf�
��7�����s���*�H�s��%i��}����`���(��I�����M��ZW��U��f'q�9���n���s̙�������QZF/�����kiKAP�/~��$�M�ݪl��؃��:-M�=�W5b���a��C`�,���є��`#�Z��{W�F����_��`i��������6�F��!�����0�2ƽ� F4�t�� �Օ�(�a �tƸ�-��n�%��$!��3���͌^D,O��9fq����
'�=�7'����N��^^��g`�	�Ewc�?Z9Jq?��Z2����OY���t��mK쭽a�C����8��52��Q����1]��Pr�nP�ݗ���0�<5�L/������}�k
��Z�)^d�E
_/貓�V��T�h��ju��8�=�}Sg��{�#TD��9�Ծ�����5MN03���@{58���HO�;�_)�݉_���b;�7�1�ܱ�*�ǓX������������7���@IϿ�/{��So��s�7!�Y�E`[i�;�L��E�?�ة|o�{������uesf�5YL�}^��ȣ������"~ޢ6#v_%7����D����|� U� ]>j�ñ78�
[f$�jMH�֛ZTނ[�!d��lS�g+o��[�{%�E&&ɡ���$`���ԽnO���¡���f�a����e0�d��%�2҅��uy�j�G��r�ch-�r�1H�Z�/��A�w\Ⱥ���f���͞K�y��\Y�}�8$Ypb�!��py�2@�~�gƭ-�����`�`9F�+��.�d~4�mơd���9?�M�R�Y4g��iP����V �\T��R��q�Gv3�A��x�vS��_(
�?)��ϴ�A==@$H��zt�dv|,ٷy�~m��ň��_�x���9��.�ہ��n�/@Ő�� H[Жq�(�z�p}¢��^�_�}\�n�Ļ/?��f�����X׻CMK�y�WD� �m�Z������X-�e���0%4Z� ��utcH�rZ>1��5�[�H�oN�4@'������50C�A���W��souxq=Ҧ���'Bx�,D��(pY,���5��������R|N\�\�l��ќ�h3!r�_g� K�,@��kAEPm�H��憣�R��W ��xں��f�%���r�S��B�K��U�
>��'@
HN��H��k_��>Q*��	�R�a[���^���:����c;�)A�)7�fU�i���� X�G��+���""���n�0�?�G��t�l�P���]� ��@LԹ�q|���a�P�ہ�|»`�<2��"y����BY� ���d� 8abBƳ	��J�3�Ʊ�l���[��f�S�k5�S�᪠���,C�TO��z�"ƒ%�W�#�U �봃 r��C�'[�uH�~���d3B���cWn���Ǡ�_�.IY�Il��
&+�k����7�L�gE�u�@��������@�8=�f�:��m��`.��(��yHo�M�9;���h�F�.�")/)� �#�` ��[a]S.t~zJ"���Q>3�p��(+��G��P��'W0̶�9�ӱ��R>�y�a���:��t�ң^�[���A�&٫����Do�*��ww.�X���0�E���3?'��Ӈ!s�Hm�tDm3���)����C�>�|��qj7HY�F�t��un/��G��0>�����"����(,��ytJ�@�Rz��j�0�P�G�Ɓk�-�Ur�f��g^���m� �.���j����8�1,f�7h��r;s�����V #��I���D!71Xx�����|9r2��r�,p�����|�a�J��tO�k3��L��Hk�c.d�����"�ۓ�9
煤�<K�H�`��Z��]9P�XXN�kT�����./���]8�m��S�݉�DW�»��ҕ�X�p�1>h~��)^t8��Zi�����,{$s+�����:t�.Q�����0��Y�c5�f��DƽL��HY'�d�~�����`���z��Bt�|�Z�<���\Y�u4%��mX�`M�7@h�E'u}�.#P:�8��*�6������9�n�����j vN�ل��d2,�����c�>ˤ��yb���LT�D#y̀٨���&�Y��IF� +�K±2�G�_Z�v�(��&�ͤ~3u�W�*�iy�v�æiǗp_uu�h:��#��jI[�`�r�����a�'��(��@�^��2U�l����qH?u2%|wx����S/SDP�#=�?v&�]�w��:K�r�$��O4�=u4�'d$2禘1��60�m�"{ˀi(��^3���������&�Q�����W�H�$�m�H-��La��}�=4�*6�f%QAt�S�SULں?���J? ��Owa��>ܹ<�(DP= A���zXWN�z��]�ԙ�0�SN��|�{��������(ه��u"���#Hn\Ό���!�k7��sM.�����A���E4���P�G��Jݍ�.;��KA�Yw�<l�����M4�����22GuǊT.�e@������fO)4�?��ab]UjQ�����x@(���1 Ș�'���7Y��� ������a��9VQ�DF���O�I�!^UV���>�n��O��p)ߢ���!�G���ܓ�ݖ�sZ��L�ңS :��k��c FWܐ}'�m��c��p��YBR�w1�n��'��42��ɛ�P�t���'���gSU�0j��*�c�������檓��lF��%!�3�O�S(��>��W�]����n��!̕Q�]!���������*�qz�^��ݰ/f6�AJ�����Oxr.��ۯYI���?U�M�w�]b��ν�=����mLE"k)ԯ��r-���i���L�X�[_���x�v�.ݸ%[�h�'�q4o.�9�4��cw~74��Qvn� �a1��O� �y�=تR\7�&Jr��3��%H�`�k�,������&����X>|^�8JY/m���r��}�D�h ���8��^�����K1�_�dh:S�i��n�9ܝ��Ҏ����1D�kɗM*��+�����P�������7���O��C�<N�:�߼q�№,K���Mbf�M�8������\��>���2Vw����SC�K�`�������4��q�Ύn�ki��&.��f��%Y���O���˲K0Řl{���ע�Mό��=����t��ʒq�i۟����Z6����l������m��um$�Ð���b�H��ԡ��]�^ap����J���:Z\�&Isg��#̳��I�}.S�L�'�=l>���ˏ�Y6a)��~�G��I��n��!���,�Q~�֊F�vV����b����'9�������a7Fz�E�S�!����o��v> mzm�^3��O��I�ms.D0߅��'�uq�C��F��mZ�K�:Ӟͯdg��or�v�]�*<��Gu?}�,^�����7{p<s
�����d�	�EZ�w#�$0G��w�I��+�3e1���U�2Lp �5�ە voen�I���~.v�_g���)�(����0m�.H����NK�@y����*�6<R�y�r6Odd�1�ZO�b;��q��-�`1xDHT�g�t�W��!�4N8��sv1�w4��w|��g�]Q��#�0��{���(�?����Py�F{�>P�DAp�,3J��iM�k�.��P�7����K_�U��ے/6	�X��If�����#s��K�?��*)�`~�|���7ƴ���UQ4�QV����@�g?*��e4�ꬹ�����=;��G����"��m�E�no��@2���= FZ���-����^�U$D\���ߖ�t��(����awD����V���[��ňO�R4=��a ��A<�9�H#�|�Ѝ���	��ٮE@h�j�z'k�+3o)C�,�}��h
'��6*�9f5�lL*�2�7�@�	*���[*�B������t��JdE{ۋ��9/xjKw�K��P��P�{|�n(�,�q�8�}'�b���� 3,"�UA�
3$m����`��$n��B��Yȏ#�}�O�7�����L�w`Z ������(c�O�� `��F��t+�t�Q�I&�^����6
�)T��Y�0�{8 �������Dm�&�x�5����L:�;4�����U�X/��J=�[{>5��ŵ�RJ[�z��})���m�9\<0��z���������.p��a�1h.�� �Q2pN�7��vs5��$H٦{=��(�J�)%�k��a�X�ˋ�7��W�/A)����*�E�mK�	x{�f`�W7�Z00�Z���?bZ�[н�t7���aB:��6;i�PZ�����o�E�7���J�t��W �t�	7���Ĝyb����\�������&���y{��5N��������% �?(���[I_�CQ�b�bW��ϰ���X�+���]:�C�ӫJ�1f�<��J����>%���w��·j�l�Jw�V��9�}�Ѡ�xb�2����y�r��N���mr��}3'�D��\fE�;�H\s�;J=����i���b�k��]�G=�#���hz�����~��c��w�����~��ޅ�E����X�c`�i�V�%()OC�� �﷓�D�T�؎ <��4�����G>�|�2���Q��FK�'�C��eb�}�!�on��8���'Y�;��o�p¡d�@����C?��H������.������-����5��3�xv��b-�~-��*��{���詭U�ˀ�ҧgNI�eٺ�WSei��CB����Il@1lH��z"<�,{=�oA>�$��ʕ��ā> y3y|́�i��<\�c�t�'�C������H5CZ^���`wU� 2Yz�ڬ�z�0��9qm�4�H���Ńq�n�߿6�P����q�����]�!�t)2m��	�'2_\��Se#�׼Ņ�hs�ς��Rv�[u����2g��18(}zxg��R��JԷ��ߔ���ۼ���=T����ߋ2:_�ܠ�����m�1y6��
�: �U2-��?�Π��z�+{��V��9m��	�lOāDA>�����r�쏻@z������A��{�p�Tw��g�Ֆ���@�g�x\"a{ �R��d�����w�3�9��H^��%���zJ�V#g��ݫL�b�l���)<�nv�ψx�Ic�������[����B�jBu*��k+���Z�-:m�ف�GG[�W�Bu�1��"�\p�p~-ï.��#�qYޮ�7����j��W�"��f�_t�Īr�Ɲ\�����Kfz����U�r}�p+��j^��Ti��Ȕ��.�h���b�ur�q<x��Qh�WL�C|\\p>�3�X#��4Z�ZK��PA�ƴy�HR����i�zE����h�9ޞ�S�[E��em�A`D�diGR�������{�Ea�ЕM�aЦ��o�!��� 5����g u�%���6[W	K����0]��%�k���?�l"J�H&*ˢI�"yƺz~��:B�aN���y��OI Z� M�Λ'7u9�hC݌E��p)Pp�m����d�ZK��h���K�2$�(0+��v.�Un���:�
�ݘ%[�ͿZ5�fB��g�����4��_��K�=7�ɳ�Q��M�.���T�ւ�x�U�b�j�<Ů���~�4��\N����mÏ1rtP����CI�p����R)�!FTX�%)�;)8څ�4�{�ّ���X�3�͓	�W?}�e����%�� �9b^�Z�na����"y/��䱑����R�nE��)9�,}��b���/H�E�Yd�kEv5ߔc;��0?`1�4!9�iz�!*��Mm�s������h��I��J���1l@�c0��)L��Y_�����:�ip�Xe���a$���1v�;j�.)C�)�M���K���N�c?�\�T�[ax����l?j�x����>�3��l�ջ]�6h6O�$����'��vN^�l)5T�{�8�7�т�'���
a`y;%�[��)�kB����,e/ՙ��H�X�,'Ct`�B[_PN�p�(����z��J�8�C��=��7�)�H:�`*C�n�t�{hE-Bp�h_W�I�*��a�n�$Z�= ƥ��l9�{�ȼHh��(�:P�9(n��2��l^\@�sS�q�R���+ y����x5r'��'�Q������#O��*3]d(�R#��nt����{�*��@J �*�)�+,�1 �&͐��:�K�Au����IGX���!���J�\����%f����:��;�Y�u=vHLqnboI��AQ5�������ӵ
��H����>���oR�51ͱ}��ʄ��Z%�bOњS�/�O�.�(�Iaa77\n�V����c$ð6���'3}�ҡ��Ȑ�	��`������L�:����L�M.��\,��kp=�iH�v����e�[��]b(Ǳ�{���z��z�E�uv���6�� ��� �*��0ÔsB;h_�i�=��ke8=�5�ݤ��)I�3��S�ݑ�@�x_K���AF/��Ϸ�Ʀ/��J�����ӽ�!���Mٛ�9�P��Z(st��B�nLY��}ac6�o�QLx_}|���`�9*�#b�U��7G2Si�㤳����s��Ĩ!1�SR�u8��IP�U]�S��w��<{��`V���
�1�����ߐa������2�k$jUI�O����»I�r5��z���?k!�"�Ɣ�y�zM��s)�E��P��y��LzLP���5���wRw4� =��l�<��ވ��f儎}��!$�4�0�uiy��I��9h_��Ы��M[w;��������s	%����a��D�&��:9NF�=|,��޾����@��`�.�jo��5�l��˼Ţ�HX�Q#��x���,K�A��=� �v(>�	��L�·>�fڎ����if��)]fb�
	�� �3���'�&�7��[������JeY��-v�����2��㩇$���k�u�6=]�ƀ^����{"��x>h�Tb(���6ț�"No�_N���N�#;9@���He�I�+f"L���������_�A9YR�fz{�Ao�~ʸ�@D�OL����sH�x�4�5�F���=K�aU�[�}S��Aʮ��e��R�d�"RΎ%_YA6��?e�/�C�aE7�D/G-��[n��Gg�1\�Y�� �}(��SgV)�$*kB�ө�L��(�Ϫ���"�{IT�B��t�����8G��%�\]�:g�@ί�5H3�_�I)zC%,Ţ�,�K|��6��}�]*�`Q7K
�@0�Y��X���?1��+;�&#�a���<T���H�P*�Ӆl�/:8>��L��j�����0VR��$���Ĝ;^J��ĕA"3ƢCX�M	TBx��^s����O� �k��FW�6H:y�QY�� �F�?�;v���z�>�q�S�K-���;+y�A�:�/;@0�����K	}w�/}���
�@�iS�eZ�ms�����q��Jp�F>3�0��m^2��A������]��=�t�O����sX����="����..H鳧�\R8��_��Tz�!F��{%�NF���q
9%�qi�&C]�L�p�?�Ф�Qb���d�5�;�QhT��6�z��\_
g׉1��8�kB�L���3������F�X�"џg�qZ����EF�!͐�2��Qd��F����L/S�U`w�v�
�7L����?-���샋�R�kz3l��GPi�K�h���jA C��{1()d�p�yD�N\/��q���WQ�yJ�_�l�� �q��jS�6��!��S��P�P�k*p��nc����+�Fu��/iJ^�����!�;�p�!�mn��\Iz��V���[t�o���E���$�a�}	I����~�L�����[����N"����LB�↍�4�T&�`������"�?������(��?:��h�fZ�i�խR��Q���A-{�z�
�*��K��$�,5��C�[�9���k�ir��G`�[��@K,�(�d����c�a��5��p�PS�����,m��U�D���b0c!~������C�*��k^B��_��t+f�w��G/�2�-�א��U@?,��"�7gxPC�2�!�]p!����u����_8��Sn
p���\�EM�Ѿ����9���M�<�U��[�E������Ds2 ֞ ~�J��Q�����5�����TgR�}�53�t9C���`ѥ�DT��;a�����}L>Z�0��Ɓ>6ƹ-����wv�r�f+���������O���;��N"<�w�>��+�oA��1M[Ǩ�dz,�/��v�h�!< �V�=*�+�������##���o:�dw#Rw,�݉0�d
��L��W���^�=O+��11���A`q]upt� �|Ǹea8䄟��]&(l �a,��������G�~�%C&�����A\�[�5���u���ϫ�Y���R�id�Q��Qm�7�s��d���L�h���\���U������*w7:��%�@�wGM1��G2	h�8�Y���V}�J�=��@��0��&ߓ 7�TM0
�%�+=ftq!��Q�������'����Y�_ƏJ���8�o�����&��룶���"g)mS�M$�ZW�d�#��� ���ڸ?Zahl^V���yH`Q��~q� �IF�ʿ�i/�vb=�݌4݈]�v�⤛<���D�zj��8U��eڿxx��zN����i��JAw%Z~��ot�C�)�<��#����b���&9tx?�,ס�0	�$�ZB�n��,��,gi���խ��L�_�G(,���N�(�)j�!�K�B9���Fgm����׳�a��V%3$���gs�o "p���oĜks͚�qq����jc�l�u��P����&�q��HSZ�M��|��k���	
���V�ge ��ϩA�h��oE<��_۪�ǡ0��S�s�i�������2�٥�ʟ�=�{�OG{�8����N���R�5��e3N��;��e3勖��ޅ�]��)>�Q"o��b=5�&^5+�9�j�{N���7����x���Ȅ�ɔ{�n,���c��/	�G;(V������J@�+\@N�f�O7�����������Ǵ/�y\�O�oA�5"@�+c[q�i�װ�H 4�a��7A�4��<�y�+<X�A��/0�1����cT̠8/�s)��+��������e@J�O�N���YZ�A�Q��3b>{H��������H.@W����e^��v~$��%�e������-����ݟ/��E���YI���>O�^�#`���*O �����d�]�����je�q����1L*�������=�w���z�	��l�;`�usu��(�$��9c���� ͤs��ԭCJ�����DQ��7����gG�ޒ�'����n�� ��&�x(9&(�F�k:n�,;�#������'Bx'�80a�[MR���=6��.�?@[9����iC��x�$�Ў*|�/�AYԉ`չ��sĳ�Jb�J����tt?� �
V��]4�-2ۮ�|�a�xO��8��
&�3�s�m��/��#�w�ak?k�F�''{�s�r�`�`:�d���O������8�<�9P��$\G~�("z���X�b���Yz���u��������\1b����차�g��A�y
��� �hK�7Y�b���,>�]�v��]7�W�:+�~]�jGt��~�8i��}/����^~�ILmR��v���A,��4��=��h��)�l[@$'8�Et�Ce L�1��+�f�NH�k�eFq\��Ey�7�� �'�ʎɢ�i���9W^�~b�@�|�XÍ��စ��j��	+��Bï�����TX`h��#� 佝I�0TX	�I�5���b���%M���54ɸ� {��7�ˮ�S&�HL��r|�����ܭ~��a9�&N���)��Y�����5Q~��H������q�k8^�A~�,�%�v�r����۫:Ö`4�=cd��e�ݦrֈ�.H�0u/�	�U�Jc��4�L���`^$	U������8xX,Ť"Ӷv��1�?�=$ߊ([R��2���I�B���=�>���V��J��!_U5�^�YJc�r������������b;D�nxhFK�'�l}=I��[�����A_�=X%��!��je�9J���In���ċ5��M���=y���ȝ�� �zi�?(�i���n�F�� �B�dOG�' �A�c����݉��K�&�*���o�[����_�R纺^�]޹�g��8<*T ��	�$?
kN΢�Gx_<�.[�h�2�(��;:��B�cr#��؎�,l~9��+�/���i'�I
�f�w(9�/)��z�4'C��hp���YC�m5m�L+��2���sh�l����!B*paiS���� }~�M4�)��s�"���j��nK�����է����Mﲍ4U��]V�� ��� :���=�"0����}Le�c���je�p{J,dp��� .��:�Z��;r��rW?���z�4�a������i
������&TO��x�۔�ꖏ���'��xM��<�pH�c[�s����x5o}��.N��C���ޫ	l�����x����m��]�aF�1��Y8R�x�����+���6�x��<F�4Uŉ�#!��7_�p�qߨ	��
7Ϫe[��,hk~�*��x{� �$�4��X*	G���P9X�G���i�^�] �cR��q%��X���VsT-��w�r`%*� ��<(ѹTGb(�t~����z_xV�
X�����B'���Z�Q�Qgo]vf��J��D����4���Of��*���K��5�a��6����N���]VT�R�����=����'�Y9	t9H��s;��������,�-�	7n ��5��kR�|�����
fS�6���O�� ���!��$:(�Ӄ$��;�5\�(�KLY�(��3�`,gå�u���ѴG��w�އ>��s{�����^���4��ji&QE�&�0���61o�<Mn�������:y_
����N�BrPO�9��+Y�1�U��QU��� V;�Z7|LK�����G�r�K��}_�G�FXN'�̻�z8<ԞQ�HސVx��<�7yp+�&�W���SB�{y�;O��:���o��o~�р'�b�o"�:��ߨ�:<k`�ED�`z����9�QLy��k��C�|w&�����=6._$�?`�O�MP�"B/[��~ ����e�c�v���{&�~
t'?��k�����cnI�ǇD'K?tk,�%i�K%��#|�����x�gqd���8@��H��6���sL����󂱽8��t��+5�J9a���Y"r\E7��I��V͑� ��B���,{"�0�30��W?�1;�?[���zL�b�M�pE-(��^1��\��΀aB�w3X\	�<�l{+{I�מ�({�ب	��y3�n?l��`k��~��7>^�P���
�~��Ӧ�I��Gڱ��2i=�<�N��څ��n�ƈ�Y;��e���C?4u������"}�/@N/�2�@��m��> �z�l����.�;��j��R�5���0!�28k�i�3���?t�h���_��0�$�ū��k�^#ө{��FF[�r�Y��ad�U��%����n><ﭞ��֏�-�|�*a~�X|�����4� �:�Pi",���(� ]e�?�A��8� �mB	�K�K��Y�v\#�m�J^�
8�&��� �@��|����¦�rL��\`���lL`h��+wA�%�]й�J3�
���o=v��੾��k���EZ��Ǹ1����R��ɿ�s����6��{���˓�R�'EW�=�;����k�	���W�H���8��E��B��tXZ�&ǓEl��S�\�ߔ���S���A��DPk�p8!6���!ʷ�;�Y���a�j�Rm�}_�|S�n�g�2`,|�6s����;�����b6�Ո�ƈ��=�aM$�$���(���&T��$b܊+�]⯷d��M�jIݗ�bg`��4E�bw��PXI�&&���xrF_�|��<+��*-g���PS"+�Kͷ�˶�ˏ	)�TǴ�꒖�t�T��J?y�[v�Px��0�s����`����-�7Y�]fb��M��'�t�rk_"Y���ЙG�պ$�������Kot�f!�� `��D�WAwJ���������_��X�j�UA�Q��d����c:��i�2��	�9��Y2��w}����1��o�mE� ���/֘J��.�ӼJ�ȵ��J�� y(�L!F��ʤ�id�+��e��x�R��#"�KnRQ����zt�+n&��d2	� k��pי�0�"]ʇퟁ:]%�l䙊�"��xn��;{|�';[�����J�ǥ�F,�q� �ή�-��N��l����6�n�x3B�g�j�/�ĳ�p������/�[�F�F����&�T��%��͸�H)z��d�6���ާ)�t���D,�(6���T�*��H�
�%��
�~,T�J\�ؑ�
ko�qX9�#_.�ڽ{�#>�r��Π�C3�R�(�!$׭3��]���Υ6Mrh,J6����:t�GSvET�����6"Y�O��{�y{�4����5��N�`M&D�����z���gP�*�+"I��z�5�lC�l��w�%X�[;�~k`�s�|�v�>� ȑ�JF)P��f�O�f���:B�J��IX�i u-�������'_��;|��� ����zj`:��S~�;&�g@@n�/�m·*�Ը�gK4��/�hU q۱�)tn\���c���&����&�G� ��g�,�
������jj�;Gc���76Lb�p�t��w��K��S/�#���I"��0ݒq�\��Y"��xFM���&,9M���&�ղ]=�n�vMR��
X�-��i�b�o5�U�
�C�������`n;��X���������#>~D�b����T��Mg��M�(��|�aN���16M�F�MZ����_OHs�Vo��ƻTaQ03��u����
�o����h�c�.<�%���-�֠��z�Ie��Z!�U����&�C�>�h�؍H��y��^`�T.B;��XuP�2^���s�3Y*�6��KRK֜`�U��oH�V0��,���i��!Ҷ!D8g�sv�:�)b#��g��5��[��L�b��ya��By��T����`e@'���B��'3W�ѶXk%N�'u�z����T/�*���Q(�06bd	^�(^w3�Y�Y��,�p�^LA��p��kZ��KX��|t	dГ�ΰ��̍'+F<���Z���(B�$E����ܠ'ӽ�;`B�����{���&����To�=(�xx�{����߬{�q$2�c�/3'�ۦ�#Bp.����6�t�LW�gRۚ�&�Ǻ���Tm	k��W*Cc���
��P��#/~��o*�m�������Jz�|����3v�B�*��T���k�����T�8e�@��,�a��S� pi�̉T������ǲ~~������Af��Ye(�U2����n;�HqBZ��-�z�"lr�C�D;,�N��-hqsDN�R_taa�$�f�=Ǚh9��rHΏ��9n��y�u�)�&���c�0��$=�s2�<b��dT��{	��g6�!�����Xc�[����7�_�(��ؒ�>
���ҟ|}j�:U��өˊ�����C�${�1���\C��n"Q��78�
`;���^��q��s���%��H
3�J�#b����a���}����]��*�,�[�����u��Cl�cX�e�~4
�D$4�W�"=���&)*�\"6١��G��i�|�Z��q#M�(�*\��/�6
F	��GI��8bH�@K`��V�Qq�����A6s���˝��i9��L݃�\�(]kzV�� j�[Z�"�%͐R�Zn-���
dW
�צ�RM�uȌ\@<�$_�ë>~��5w�Ni�/�� B�U�e�����2�d��g�t��8�'zD���j�QP�D4�gfBf�/K��+&
E�ک�]��.e�uI��l;fe�~w�`au������=�u���!��b�dfBV�(R��ZO;�a!��7���E�l<a�ɍ�T&bM��"��༴Χ�?c@{��^N.�Xd!�2
7e1�����4��X�����K�r�'�$�Ȕ��V�a��Xw�)�9,ڐ���Ժ�+U��G�;	c�.y���t!�׺�j6�)}�������d���^i^��A���u���h�l�g����z�u���ڹMw�P��^�#��d�ԏ���h|���2��z!���h7��v�������D�[��&}̐pSC��k9�RS�G��
�^��ⱆ6����5$*l��*=���a�u������'��@����Wi�˩�P�:��]4��.�I3d�`�uyu-���!a菹��N��rn@w�۰���֌�)x�Zp����:]/�_�a0#�۽�4��qZ�@��]6�z՝M��G}�	Dj)/���O̙A��M���0�V}9o�LࡽJ���^�𓝌=1eAh��ϋw�j��t+W��	Ҋa�;��][	���a4�S�������g|�ݘ;+�ٴQq7�������� qT<���(�Yږ���L*�	Ʊҡ"�����[�g"��7�?d	V����E�V�=9'�����d)a� ���5pb��F/�n3 ̹��WAج�`��Xv�o*
0�WAg��䉘\�Z;ʘ��.���n[�B����� N�۩�팝1(� 8:�3R z`N'2Oew��s��� ���^��	n�Tݕ�2} ��J���ݮޭ���})D�vJ��d�h��7�Cju�n��+�����a�R�V	��)�?�^�y*������3̩�ٮ,�qp '>�����sC,�ʒ����38�`�S����{<�/��I�|��q�����}D�K&{x��n�
��S�̈j�߯���Ǿ�� AЈ�{ #���j�H�w���4�J�/A�Y��ݗ#��c�@���6^���H�䚽�5:6�Hv'uS�iFL��.��L0�^�r���`V�M� ���u�H�(!,�B-��GQTH#d�<%Ng��k�r\��b�*S�zky�����fxe����_�%bڶ_�����/Ű�ւm���PƱ^���2.�ف� ��b�+1��ZX��̼eȱT�Eu����9���Z�$��n�拙�V!T	�IO+�|)Ђ�!$yk;tS6LD�W%�~����n��Lg@[H��~l��{��5��,ݗ����%����
��ٻ�bşnX.}�O�M.�r�I&���Է-=L�:��W�A��gZ@q�$O�[1o�����-Pן�\��7<ǙBZ�2w�\%P��F��K�:�nh[�F���GѾ���/va����rV���O��8(��_ca����[Տ���L/lxpK�/ẕ���(��ƪ����ny����-査���4�Q��&�^r*F5P�M�P���X+j�:�M:ȉ�Ux077�~�>1�s��X�1 /��8;��>�G��4�P׎ �3qvK��1�)�L�u.���ϝ&����&�#sM�����=��vl�z��>]�cU#�&�AKLw�2ڑV5 f�e7aO� Lx�G%9+e�����a-�R���
���ۘS�ز�1��qI럲����K?;�ۻ}4��,�C�;
tX=KTE�����M��$���՚dx��SP�Q H�j<�jH����LS���O���Q/������W�rE�
�dk�l ����Q><0������+&OI6���3�zB�\��c��,V.���R=FH������	H��*t�e�(���;�:2FG�Z{d���~)��4�q�U��S��f�{�2�p���)�����Mh̡r����@m��*��\��m#n2m�cN���.��ۨ}f-���M|�8Fu[��+,3��U-��o��t���յ�G6�!�D�@�( ҉�ֺ픐](��:^>�b�w����M��e;���J��dr�L�$��,��K�����Q��#j�k�[�vܻ�E`�v�7:�>�M����;6�t�(����B<Ě�Я����ۏ7���!D��{'2-#AQ�a7�A�a�����2g��ު��>�0��_6��a�p>��i˛�%�Nk�g�HH�yq�5���Y�������f�zm�uU���y����(��S+r���H ��=���~
e!��䑆���"��1[��n�{��M�,��y՜-d$7��b�.�c���%�OZ"Y��F���P��_P~Ѓ�d�MF�(Iv�}��=s���q"�N�-�b���3����w�5����]��u""Eu�L����g�l+	¨��1�㉑Lv�r�ϟs)�㰕C��1o��V�8�`V�&$�cRvX�%��A�����X��J�K�=��	 �:�Ɗ`����&2�I�2�1Av~2C��G�|#o�Awŀ.���z��/�5�q9Y�x��Ҍٱ�{Kd����v����UT����|WbSőYX^��y'n����m#/j�,e�|�6�)��E_sh-�Y�4;�8��۠v���ٹg�cYVy��$Phx�>hs���ʉ	�� b}������v�xg�����*��S<��4�Gx�\�)Qѹ��B� �U�O5�Q'��.F�.Y�u�Rw�K�RZ�1����oGEjX]H�d^4����
1��Z,1dHm.L'��ʐ���_��JsK�@�IBF�Yf3 :�� q֏tcX���7A��1����a�p��
 �&��|)��}�WeoU��|6���÷�2��ZT"�g��Ir����u��c)llXu�6��d.����hw[�n	���p�Oِ�I���E�P��V�,���oD��iz������q"��Xr��;Ŏ$?{q��t1ly�&�4z�E�Èpe2'/�3��5�O�3�5<�">c�����k�$���,�����}��
Ҍ�S�2@��,�^w��FAZج I^�[��8���cX�/dЖ<z�\t�m%>|�h�Y�$ܢsܘ_�۲�s�8�i��R�<�)�z
4M���������qQժ�s���B�H��GV&ޤ��q� �l㋊�4����|��ǁ���2��OL2�Yh���ɇ+l���b=��%�:��G2�ic8�k3>Ϙ�w<iH_�t8�%rCy�3�/��)��Έ�޵�:��fD��H�$*^=�:��W�E��7���W����_����ϓ������8}��i�?��,�����U��O��iwd�P*�E��MO�����6��%f��ɶH.��*�|�n�רX�+/�a�ӣ�_�|�3�P�P��"����ϭ7۵Í�G��<�Ŝ�ud��Ohk���������hgͭF��x�!�wK��N�S�*8��	6σE��,ig���5	 i���r�� ��{�)��Ν�a}�I�攓%��b D����_X(�D�iD��r!����6�R���S9�:����	�
��ȩ�p�n�I�K�!���D�[�#K��)Zy���	dh��,��n��.�xn�7q��\�6�J�+;�E�c�[�ۻ�6Qڿ
Y��l��u��xrө�?�����Tn��~y���o�b������������b��־f�eQn����^��'b�lz�ZDҟӝ[��X� \}��eo�h"P"]LebkrT�c��d�"j�U�~��t���$V��OM��Y�r��I��,�&�p2�f�) E��J}��9>M`����|�|����.jִ|�)r�L8k�R�0}��2!�p;�n~-��Ԃ:���7J���_Z�ѻZ�9�{�����dUy�. ���}3e��Ro����b�G�0��ǰ���?hbB:�0�	�[_��/4��)w��^�(�3w����C\�iv�[���R���r�/���
�N_*_���D�e*���uE�Ь@�av�uO���N�i�夤��4���� �;ůq�g��][ޒ�
viF������^�\�Lyevxɖ�phVּOҜR���Rߊ%T�	e�a�������W�]~V/���M�>�Ñى�I��,��/�q۾p�EWρ{����mz��ru��Bs�q���ޠ�LFV7�Ri����3"Va}����LLI<�Sv�3l�G6�k�k�_�6���n#�Ā��jF���6a
dd�y-�Bˑ��q㓈�H��G��+r�����,9{�λ��GS�p=�[q+c�㖲i@���r���*�����+ҥKI�_��=P4���_�1k�� %�$x��� >h*$O{j�{�b����������7����c�r��[!�h�-w�vE�O%�"��{��|�o��M�S���z"�-#���֭�Z����*��13$��GhV� ��|�9)��D2Y��iІ#L29i����w�d��G�%��T`�L4h�i�0AZF�}��^I^s�o��i��Q3����J]�ҳ�U��v�c��U�v�5]�4$0���j!縂�$|���E]z~�B�$90���n�����f�'�)�����]m"��:#*��:Ơ��CEO
�LK��P�
�:�X8��`f<�Dl�+���H��|��Ϥ�#c�yZ�}.�m)�Gj|/
��l���Qx�d
�H+�W��Jns�p�t�@�����KC]�8ƃ�xP��á�uָ�5��D��CPETA���n�8�/^���Z�ȿ�f����[�<��W����.燰r�^}-q	�#���l�s��ͧi����J#�/[[ �7��Z� ���O���H`��Fw5��|�{��,��򏦠��:�Ra� �
��p#��%��\:�
A5:�_�|,�>S���E�v�( �|7�؍O��ψ-i�e{!ӌR�])�8b��-��e�	M�L��z��[��Jgz_-���FC�N��ݗD�l_e�S߇����n�����SF�#��[r��d�Wh����7����m(U��;7@��[�����ް�����ٻ@ix�1����f�"nؼ��u�O�Jp)1�+�Z�&KL��?��=�P2��ʬE�9���ƀ�:}�]����?�1Ȅ���ܬ��^4р���/c��nv�[
	˛���H�SC�k����ҍ��+MTg>�[~u�R�Ϯϰ����)oޣ�/�R�xZ"�9ʣ���>��8��cIOX����*?���]���2}p��	ڍ�V�"��T�cDIIX�	��"��Do��Q��Y�[���2��<�94���IqPcMdDXrS<�=3N$���SB����U�Ӑ�>��<1���b�T9O���&H
1�3���ʽB�_�#w�Y����(OJ�#���*C�ʖ<צ<;b��6gD�+�@��B6Rzu���p$eXd�6~ֆ2ws=��c�5�FVR��H�rO��;�h��:p�Ao����L,%�4~u!�#7��O,�rW����{�fYO =�I���-�ݻ�S�]�n�3��o&0��2B�9y�N��:_?�dAn�g�P1����hA%h��
"�W�����r.yR����s_�joI�i���O�:-^W�t�bR�=�\!��m|�F-	˞y���:�Цփ���ƈK3��E?"����0Qa�'�v됝*�	�I1���K"�@��r�i�@a)��g�-�6��Eg�H��|.�
�l<��čPᄽS�S�����<�X�f�̀^�@�{�M �=cۉ��b�Al�Y�űEF����ϸ���aF���&�
k��t��FʯXtdd�)Ҕ}>����30-�ʬr`-{���\
w�@M���J9H�'9ܥb-��xfƟ��ڗOr>9�6��<D��8h}�mGkV�SF?����#1���T`Te�t�����:�	�g.�I4 9Kzz� !zQ ���ء�K�A����H���.§�޵D�[a�S�E��k����ּj*L�4�g�S�
�VDV'?@fl��9^�JB%��i���g/j��s���*Z���C�M���S�����Tߨ3�ę�eG}� ����$�gL�;~f2�4���+�U2d;�����Pp�c��Hh����"el�+d�-����w.z�f��ݱW�]�֐��I�4�OI6�>6u���&G(�@|p^���/�Y�qKQ���kB��Pb�B�������$f�/�\� *��k�9�]l. �H���~$la_ӑ���* r-9�g(�^bN�ZS�t3�O0��!��QE"A�I�L wv��)�� ��?t9�V[��
��6~�ZS�3(8+�dz�f'4�� ��h�(R�,,��Fsuc�]칿�|���~�S�:YɣCj�h/XX��Ju)� 
�����: �:�����<��;�
� C�[�А�;-6�F�T�J���R�����/�3�N���^惐J�$�ίW���ipL�Ŕ'� ��ʫba�Я4����|U����Cx����oh��b\X���
/	��K�N�Q8G.U�Q�Z�v�e��h�FB�q���A�%|C)��ZW�)�ics�v~-����C��;ŝ�H��"���/�C��v�!�j�X�v��1��,����\��~����a�L�N�^b>�h���L`���2{KW�8�/o�zŋ"�����+q� 79��nO��Z�κ63=E�T �(�\R/RI��6U�`��ڀ3��k:���g��@������x���- k.��;�{��߁��5~���kػ�L$�������ϣ��(�����A��D�)Il��9@�	����.�b���u�>ySH�秈I�n4�9��mjG���
�L.?s8H �\#�i�-Z*Psa��Ar"x�������[�8��/���>z������(�i�he�g�MƑU�\W
��� +kW�ٴ�0:CIR����'���FU��w3��l]�	��Jr��b�kr�7�~�ѽ�g�4�#<���6?�0�y� o��)0��J�۾ɨ��Lc�شr���}H7��Sj3�'�ҁ�fْ�-�@�gW@�ҏ�4D'
�\��^�!L��(wiO�D�ی��z��v7�g��0��*WOA����)����&��E�8��>Iޯ�}rQ	��ԟ��-����su�1Ȟ����cp��mU<�����hc��3�7!��"�s�aZ1B���Ge�Ts|m�?��#��k�%A��z�y��
��h�DG�x�T�s�[��*%�Pm�Z�vC5P�^��ؑ�՝7���!�k��f� [b��I�z�2���u��ك���$���Ka�p���[{��2&��9r������%]3�����9ia؄1;g���0�h��L��^�W��!0Ϳ��a6���>66�D�&&��)s��UdcS�PO�g�O�IYM�{5���f	���'�ۊ�?��2�6��q���v�ᐁr��۱mA��R�rńj��^f^8&�P/�ٟЪY�b !<xq��ë@*���U�y;�^h(��A�ݝ%^~�2� %1&Mj�K�khن�{$��OwFޝ��Ś-v<T�3�,������=��/�v�_���(S�,�$�9�>�^���|���Ŗ,�(��7�0ù�%cF��U`�V�w���<4k`~���~ ��=ڬva���n�-/�v���6�����V����Gƪ���`�8A���H5��ҵڱȇ�4��k<��IbȪ�a�9�o�.��r�5�c �|�]�Vj�?#�Nh���xUA�3��NF���,r\�:WT�W���9�Y���fX�$"cs����Д4�\�6�!R�v�r��ޚA��g�# �%��{����R�y�4��Z�j�.����X5�Ҩ��${Ӳ�3�BBu�R{��MHrHDfov�t�Q�L�ϋ"�*[k����JS�C0m�Z���߶�~�/j=�ϧ��O�*��H�mr�d	~,1���G�Kw���;)��F
��؂���KP5�(�,ϒ�I~Iz`q��,��ka��E�/:��S��L�1��6dx���F�W��Q��1��}~9�nk/i�j�"#�l,87�7�QH3��~��n�$�n} ����(H��tҁQKC��������f-
��zX���)�#G�Y������I�O8\�����7���mT�ˇ؃S�5I��	�
Y��$١c�l-п9�[d,��}�w?s:��T����AL=��2�wX#����Xz�J_�"�FƭOa�X��Q(��{�c��h槏
wz�r�іdVDp��p%�9���_�����.}_�Ѧ�Ǫʤx�G(� ����d��* �mi�,f`�g����4����ij��;�z���)�b*F@=ɬ��K:���!��lӤP[��	���)�)�T��{���n�g�'�*�&��N�� `.}g�!�,(�����o�����/�U��΢�����Ҽ6i�$)?�q~�kP�y\�/�9�ԜC����}��__�cB����S�E4�]R�?<$�~�Lx�hE_�3�P5l��$���3�1������fgX�{N3��1�v���Kañ��ĩ�L��:~ԃ\2�H���K*�|�<.v��>J"0:������=��C%7��Ia�/߇~k7�4^!�j�3�zp� ��N���5�vw��ۻ�'G�e���P����me|m�vy����|�}���,�7z�#;�VY���-�����^���NI 3,��S^��1̭�v�}�N?P�kW3���i�f(�s��%ɿ)+���!E|<o��;X�c*���D��_���r�����>�����5�OT�7��1��\n�6"��:f�p���熄���.��icM���Ǻ����,�%�i�!|�M/4���VG +^��7��B��7�r��Άgilc�*������nh2��S���_��/��nh�I�<kC�-�$�C�kCh�,�u�.v_n��5J��I� ��C��Zi�[N���_.;8*w��im]�U���b4����|�Wr���f2�rt����OHXIye��>��C-l�~�:�qM���*^3؞�at���S�Z���f�A�������Do����2J�!�j�"p�_b�U��N��O ҟFI�	�l��~�ʎ�c��c�棌����W�ݞ�����"����6�8C:����c+F����*�u7�&J�v��ݧ2#P�S������+�0�I`P��Hz���-�e���ş����e�߻�rȗ;��a4lat�\D�O��\�F�N~rA�#*�׹���#Y�fr:1�����W�4�^����J�h�<S�bt�M:!rNa�t�8�| ��@���N�"�1�Œq�����-����*��8���z:;k)�&�����g^FD�h�y g�@ҰԦA�j���22M��&�s�e������J���'A̸�3�U�����C���?gy�x.�7������8��s��0���-��6Y�r��5�߹8�Ħ�������f���;ɜ""ի��o�\��<�^8��r�.a���+ �~���z�!f�_�e��יe�2��Ie�
����l�* ���d���)��Ua�mAu8�iFAg��{4�wil�G�΅��p�(�=�e��Y1�AٟZ��:_����q���ǠG����v���7L��(�K��ϓ����W@���6Ң&Ak͸`�榏#c� ��q(����|���y�m�E�cN�;�u=�A��/���|����銷C����S�v�k-)�'x������);�pd!����" n#���\��a���s�ʘ�| pnj��S'=Q�H٫T���'ɑQ���]��`� �(Z��ʏx`$���V_��^�����?��J!�U3���6�j�d�q`)a7O��e�!�O����� ���FLp�c�c�!#�����ANY]|�	��7|���s���Z�ln����b��t�mR��%�X]9.�����H��'R���ˡ43!�?�M�1�i$���K�QID��`��r�.�Clt�i����<����YS�F>�Am��/b���dn,U��@�����[4t�8���m����Ր��=l��[�K�8���@���4�zX�Ջ �ּ�wi�S�*���p~�����d���wy��WC�Ɇ��l��A i�`A橨lǐ�,��=Vm�?�C���}����PCO��W�хab��I[�ظF�U�J9��05c��h�g����f�*�,�|���Aǭڀ�f�9��n4VS�C�+�#�l��j�*Y"�1t�9�|u+��+Ś��o���u��j����|uL�6iK�d����`��7ϫ_u�h
�%�[
It�Y�M�bTN^-�,-�V1�tE꤉��h��g	���,XCSe`��b����e3�b��0��^��*�@W�m����Hd�wnZ�t:�f�
��v����Y�sڰG�z}V�.
����E�Ns�W��3����+��^$T�ES'l�axZV��{:�X$�}�]@�z��[x3�n��$���
c�(��H4���k:y��_*�"n�G.[뤅ݯq�A	���>��/�P@����x7��`@�@>	�N]&�M�r����,��o�dE��t���o��ep�@rS�J.Ƅ&�3�}�0Դ.�ji93w�^���%	J��pN��n�EK0��B(�I�~9����_�R) ���Coj���{��7i��7/�����}s	�$G����щ'%`��f?���,z��D��Tj�Ѡ^�?�\�M}��S��^�?��B�t�����j��Z��w�w�OҬ��S��Fk"���0��Z-�83�t�p0VvD�a�%c���`oL�:�lɧ#��吚s��.��_j`�׭�%���)�"�X���&S�yyDoQ|s�3�_T��V-~d~N~�F�U�";��v�2�'m�+�AΈ��;�:���Dr�[����M�W�W���F��V�=�|�V�J;c2�
vg5������5>�x�����aQ}% ���l5�w�ۥ{�[�\�+!���<_p#5�Rx|�UjeҮ���ags�o����Z�9p�U��)���OQi������ްf�0!|�ϲ��CZy�'�b@\
��^�P��t���}�s���@�fX������Fl�-p%���]dI������c���B�ڰ}�f��OcԨ
ж�p�nn7��px[� A�U
��P1�-�}�~r�e�0�<���ƻ9|���QDӀQ� u��@�C40S�,��1�)�3\ܳ�灇qkO���W%�\c�qS����L���!��&��a�$I@i���ϝ�����>"�d!r�u��r�=���\��P����F��z(�C'���֪��L�`)7Eo8�.?L&b6"=�QEe:�0ǐ����-!�}��D����� ��|�N�m$+�8t�$/؜rZ���R\��b���ߺ���7�OM�#�Z�����]r�@���@$v�ݘ���+�Z���&���7�1���_����BvS���΄,nΞjW�E>ۼ����,q�Ҽ��-P�'A��a��|��kZ/��]AJ{3�p��IF��v@�>�bQ�p����zO��V^^���h�ѮFsѫ�K���rf�,B�m��ŭ��@�"��̍�`��|�v�x�g0���4�es
.�o�X��l���/���.L����s6��/�`�b�Py��=�3}r�Y&���Cq�w"��i�
j�Փ�F� ��9
X]��(ѣR�����4V��of�+�N�ڸi_v��Y�a�ɀ�o��GO��ւ�$l�`�y#"�J�Cw�&��+��Dި˜	��{&4!<��ن0�;���r��GG�t�.��u9K�He��e/���quW�d��%��T�	_��:-�AD��u�YY��f�FD'j� ��F��S��e���U=e4�{�{6�$2jR��o�W◒?)���Y�R��L��N�n�uz�Q8�s�d���P5�	�m1Ű��tJC�I��M��8l�RFڌ�����ޛj'&�Z�6 9�4W�_��WezT��N?c�%F��W��K�a*��6-�W�R��+բx����7���������&��C��|���o[�A.�T���[�-��鏳d�<e���	6E\�_��!��[t}?��>�z���u|�#%�Z9���<*�]NV|�i�d1@��:X��k'�@};
�/{����
'�u�=8���(���a��SLi�d!GN=L�/�QX�v�V�@�B<�Sa�YC�F�|7i4�鷌v�w�\��q1�P#%C���y��q�Y����_�6\��yh]�#m�������F{,���F�`�\c�O��~�D\U.8���kHO��O܏5�e��{���5�
��%B\�Pd�ex�g���	ٛ%>Q�tm-�%q�oS�Y^	穊�L ?{��R��n��,&���X5�V{�_)u�3\�����Tmx��I�I�7�C�.�J�w4�1x�m$�r�&�C��q�F����*OVE"��P1Rs�<�k��#ₚ�R`�Њ)w�v`%��7~2]o��Ԕf �V�!1�eɌ��
����1#	_U}B
4P$nZ�����r���6ZX4�q�%�b�"�����N�h�WwYR��S��-��`Ү}0�D�(�����)��mʎe�}�B���`���#���)���I/��<�1��_��%��X=�s�D
��b:�܄��R�Y��Fh-�p���C�M��@Z:�dћJ�(KF01&�zYkնaC� �,�V���T���{���m����E�Pr�rd�1|ts��}��ƏV�ņ��Ɇ�U��X�wq�� �mw��U�6w������S̭痨��֑��{Đ��̿ߌ���bY���z����x�@�UR\��V�ɂ�vGR���ؚ $�/��F��`)���:�Bl���(*1M8�|��լo$�3���Mliӂ�~_���,3��$�1���brV�[���V�Ӝa ���	q]����!�Vn��_1�[��ȋ�N��*���B��d�ː��ާ��=HC�}L.�߯����tD*�]���N�2���A�-��y/���i	N���;M�u�guYL��t*���`[�Zj�Ac~�o����gq�8�>����vASۃ�e&��/w�yxi�r�&���QN������gR]�H��+LppR!�oq5�r�{�7�\��?cT!��D��b��S3=Qf]:;U���G:�l�y��C_ͽ�o�>����c�LfY�$��̤��.�9a_��-�Ⱥ�$��zم�֛�~�C��LX�K��今������ସ�dP���T������ m���vU]�.�{EB^h�Ms�>�Ž�g�Ь���k�I�|M���te��O�"+S���1c_�a��txvd��N$J:M=���j��m��X����\T�$��g7�]���pU�{RAP��|� Λ��	�k��G=����-{�ǖuӡu5�SW�b���9:�l�%Wk�"��Q���4z�U��$&�-])p���w�����;ٟ1�*�; ���<���|O��A��9X���!�<��py�C�רMO���xH���ͬ��t�h�}ՠ^�.v�׍m�vx5����`x��T�n*���o�#p-��jN�&�Q12o/�m���az���˟'��:%���G�����c�����ه� {�Bރ<ݱ�QTv��S̫5��T�!� �����,��E�MLxZ�b�
�YB[���L]>v�c��W�u�f���-�W��Kb�8��ʒs���:yO$��k����2Yʌ�Y3b���?A;~:(�D&��
L?5y�����q����L�_�v��8B|�Z�ع�^a
|m���V[����3�qzG.㘁suB`�Wg�!������
��w4�/�[8^.��ֆ請I��f��R�[b=!X�.|��Dz��]!F���3�?#aC6��|���W�aI�~���\L���֌�`�o������ź�b�>�u�)�y�'� a���Ņ��OF�0�m�f����i�xG�A��:�L�?�B����:Fxf�N�i���Xt�T��u#՞ۏ\��n�-:��w���3GDR<�_R.hɴ����!�S0�V�gf��#�	K���-�n:�rV�<g/^���t]��(`�|�LY�!�/�h���8ݤ�8�`��3V��n�`<5��0C�*>�G4�Df1����EŽt'�ů	9o5������� �_���Y?5L�
���%�p��w���2ت����[�^��GIp���)~�F���b�M1��Pnb�-�lN��e��r�T�\�C<WO�0Q��^������N���3���@Ãs�i���ބ;���W���k�G���)ĸ�g1 X5|'h_/]t =�5�.h��J���T_g�M��f������?��Š8�'*PT�΁?�[��!�ςؐ��ȡ�̨�ޑ+�$*�Lk�����y`�N�GV�j/��h���Y
�8Fb3n�U�5���æ�C}�̤����b!+���v!C��2�T��i2^���zDI�{\b�5�K����ny~`�k��i�<���Xޝl��{�� ʻ��k�� ��� �zl4<*�����$�+�gRv�pWF�� �_v )V�g��M��NoS����� [2��sK��P�+������$ �:|9�T��Ҳ�J��_����Wa���N������y�@T\��|!yl�^��r��Ǯ�*|���D��I\\����渔^�2�aĻh~2㉡K�R�0�XE��#Z�_/R2��&�UI��
�6�	��������:5�G�ᝰl5�.��^��<9�P<�>�.:@���q�F.8��%��u�k���H�S0�>Ri��e��@�`�+���w��4C4/s��)B'^��ȧ�.k{4�'Ȕin2�#�v�P�h�|�f����_Vd,�'�Ew��� ����Vt���?xj[7n�S%����8��/��f0ZaZ�TSi��������p|�+&�D�0�>��@��r��6)'���g������{�ڍ�$�zt�����c������ܳtMH��O�������d��1�"���Ҵ�S�b��x�gJܿH3����hSk�Z�t�� )@��s����ß-�'���&��7aP��A �~q���/lgg��{��́�8�R,�F9N[�0�Ծn]��x��٣c��z���٠\�^�1v��Y'� �7����<�x����4�h� �͹VE,؉��0$��L���h���>���@���@�w,���m,Ѵ��P04u�`��0�\��	\.�`�֔E�E!:���Np���'�Ms�������YJ.�.��mmE�۽���,ޓx�!�գ��6`<w������X���bOU���p�\ԍ�ZY8���ى;�$j�����2��-���CO����F�t���e��z���?� ��
n�ŧ�!3c���;�,�ޫ�f�O1���,&�0����Ý*Q��$��Sڙw@��R;�r@�+m~�r��t�&�Wp�茙l����҅x䉽f��4=�I�Y�ź��5C�����ŷ��Xk�˴��l=6��7��[!�<���.Ulq��?^�M ��85P��Х(�e��Ot���uΚx�����Nݜ��n�_L�PP�ޅ@R�%=8v^�X���,��_慬���1�Fj��=��r��P�j��U�������J�y;�;#j�X=	X@��*�0`NFߖШ=�i��<��f4��B����m�^?RR���G�O &	�cE�{�*VLC1z/������rǘ��T� z�
���l%(	ED���r� lQ<ь݋���V�P/�Az�G�V9��z4hr�|�ìw�K�T�[Gi��> w�叇.�JG�ɉ#.�,׎�i�O\J7��aAy����bV�N(��خd�����8�#� �j���#A���tӈA�8 p��g'⊵�y+�n(ۘ�����{d1W8�[�8�Q�6��S��I7,�8a���/�^�����q,���O�>���Kh!S��.�js���C�4f�S���0�I%·�<��p�I��Ӳ�C�r-{�9B�����}�D�u*�!�q'd�1��0l�x�����p�i�7�],��
߹j��K���X���j��Ɔ�k��l!C�3�o�r��c�\Z�$����d�����������x������OU���8�m�j�Ы /8�cZ�����0�Q�i���Ė��=D�j}&^[^�)���O��Ks
�A�x(4�5v��u��6E݌Me��
���Z��OmV�Z�����˄.<��l(88u� z:�Xy>�?'a�ؕ�]i��/!����+���@9���{��6�5M�?��!��� �P�$���W_'������`����CдЕNQ����q0�/G�R|<�e�^Ā|�O��r�Y�3�-*����#)FR�g&�(xP����97�I!�G�/���,���e�|6�<�����E�9�d�*��]j�kJ��c��'�y�%e
� ���2�T��u~n`L�HS���%�Fe� r	/N�f�w�ƁR��/������d��	V|Y_Jsb?��!:uѝ�@ ~ܝA5����ߘތ�����7	�u��}E=]=�wVu�k}Q+!����iZϖ� *�#r�.|� �O~�U�"����MD������HX�͍�ڸ1!)�6)� ����� ��l�"A�Bu;���5�4�������(�K�z������)�
Qw�,m��r�W ����u����@�vGCj�J����LIOO$��4��e���Vi��?�䰷�e����5�MՍ��*hq�$Z<�T7�w�-��3���"�"�C<�z�N*��f^��ųV�� @��b���90�nu#�[ϵ��'�^#~�ЉA( ��Z�r�s���g�<�9y$? �Z]�#>|��hf��re�F��7:��![4)������@��i�_�[��&��&���B1�[�����}����(�m��Ⱥ<~�#��RBy�ټ@G�h��y9�|�4�&��=��ۉpV������;3 ���wW2v�2b��pju�Y5>��H􋫉�E����]�6*p������g���`fɓ�k�O��_��/}R��1]�9^�Ǚ[������r��I*��O���m��s�����l�c�r�nM|��V�o�i���|e��Je,Ř�]�[u�{|/;7�&᫪]�э�U�b�χ���J���)8��D�����[ը���z�N�[>�B����ŗ�N�g�Cv���>�i�|Gku���^i��E �L��;��\2��l��>�]�6k���/��+b�� ,�ݷƩf<Aű�7]b������&���%�2�ۻ2�0A��rt;�N6��yԩ��P|�N�AJp�^�Х(S� N��F"��vM��gd���'�Wb�t�y��|�5o��Q�O��́<�믈�`��D��;�3��o6�^�i�����z�Q�~N�I���pvH>7�?�x4�0,�\h��
-5w���B��B��O�uF�>&�#�+X�R�C�݃qh�8������A]��3�fp�ן���gک���u�)an�m2�=�Uo2����,�������U��F����kpS��8	��$}� ��j_�,)����#��vl�+�*7�%/�<D!� ef����\JY�Rp<�ЋSa��[��ֵ��ދ#��)7���']�\�*��Z�5�6́�^Ѱ}q��Y��A�쵦Fc��ܢylg0?!aAy�����y#+�4�Ύ��oA_"��r�*l�C�m��]��ʪk**%�-N$K�:Ov6�.}�Qo�!}��A�����L�M[~�_���G=Q�g��l[�B�(��g
�g����B[�&�ϿM��	���_�E$�p���f�-1#��6��^g
J��슛�9�5	]�f"����.��������K#�ސ�L��"5u>JyB�X�Ǯ<����2�}W�^"��K��t��$
��p��O�qi�9U��h+V�	]%Z��DHB��ǆ܂��:m�'����1 x��~���:�sj�組�<��G!#���n�� ���o:��.���g[��I��u �װ��\b u2�wMc,�}�4�:E��y����jA�8��&�Q�8+�0Wr�1=��5����_��=v�:��ʰ��VU�/!�⢧�TA	X�P�U�鸽�R��Y���O�ZQ���I���?a�?[c��<:xPXm�?�W0.Z�
̢�E����'�02Z�����(�� M�??��7��R��%�`���������5��hQ��._	�VJe��
*e*��i�
�}�􅚊6�M<j�'7��S`u�z5.%��@��k"$,<)k����ltb�� &|��x+jS�3tn�A����5o<�p�^u��ȭdG�]������y3�s@5�O�ezb<9\�
U��`X\�K�h=����+7x��<���tPW��l�fTt��-d;�O�?4G���)��9�"���t���0��y��c�I�>I܆�y��H��a��1�����U�b�3Ua��:]t�1�OB�-�����WF�ʣ ���<�����P�;};#��7��F�n�E*��9`�^^������]>o�K^w�Im=�=g�m& &S���n��ƀ�J��,�j�_��2YHy��R��_��{j����<X#]���3�'�6y�Ȧ��m�7�t� >6�~�`����N.Ưh��A@?��O����z���4�L ��f������4S}n��O|����q�ל�|0�䔹8X�P�;���"S\m���^,��=Q2��pg��N�ɪ�&,L<�+·7�_@l����/E��s7.�'}��Ze�b`��ǣ����5��	@��G���T�8�LUV]�k?����-��hk<��y��(�b�JD�tS��\�#��}$�ۘiWI�b��/S�̆�)��LP:H{3>��`7zC��+V��~V��c�U���ի�,��5~��0�ٮ�3��N�����w$��}�0<B���!TY
�A�)j�������#�N�^���?��:}��= ߓ�����K�M����cL���h �����mp�$Pb���2��� ��A�S'P&�͎0P+��zL?)\��͌�C����jRR��frĜ|vx������w� �v  �l6J*o��	��`ɾ�lѦH���2�\8�b�"!,�����}$FoӪ戳쁣� ��g�"�@��������"H+��B�ͳa�%�����x���������:o�Wy���&h���6�w�dTi��3{3#N����k�a0C����G%����G��,��X{MxD��u��͗(���!L��`��{�a?����+���Ig�q���BV�o�b�x��O�(XB��` ��*s<D2���� /��6nx��%M�ď ����7_��7�'��6m�JG��<6DUr�����	���,�\&+\�!�$t~����/�]4$W��8R�JZ��m���l}�& ?�w��jVKxM���Kd���G��1�:yO������J�oO��?|1Fxizc.�G�5iq���Q���GS�
�X(��6��l�SQ�>�,->(+�<�턞y`���� �Vo�jsZeƆ����Ћ��-�hGT�����?�,�*�����5�q���5���I9�ഖŻW��/r׫�v:�u�g�M%
N�d|���bע~4E���0�ԧN�S-���hI��C���k��$�)�Fkԙ���ѝU*&9���u8Z��P� ��[D�vΓu �{D]���%�Q{�O���o�`�tQv�S�%�F�t"��L8hG�w���ׁ@d��)��%����Ox`x�_۰�ԾK�\mႨ���dҮhPl
��i4c�͌#�3sƘ_��G[���-0����\����Q����G�oO�+
J%��wEE�OQN�$��HQ	�>��](�1� ��ʓ�2��q|ld�.]�j�aP�/ʑ�*i��i���c�=���Ln�@ ^޼uDެ[��H�ў�0�3U�s+�㆙9������P˕�8��A���歜*�����ռ��Է��F!	�	=ͯ��U��!\��&g�q��S������}h�B d�M�2�ZW��t�5�Ѿ�G���{X�ÿ�3)Wש����1��!��i�&�Js�GϧRƈ	`��6�%3c4/�-4��rJ�D�����c`�&�%�7�ak��4��x�(l0i�\�x͢��W!�J�A���t}�����/�k˴�L>��4�b�Ș�9'�Ȼ��D/r�44���
X�n�Px��Pvr�����<��O���Ÿ��pJ����̠2����sd&h��ؓطF�%�X���[�բ�c���(+	.���!c%���/ʦ�9[��0��4�š�d�FUU/���YZ�R։I��a�/�D�9O�b����������� �v7cѵ\��O6�o��ٳ.��k��OXpk ��x����5�'�
U����Rnʈ�2�JׄT�
����0�qEQ�]�͠�c��� � ���|Gf�l���	X�K��p!d�Lu5Z�<���nxl"��Op�d�	�q[Y�ߨ��/�>�<*��=;��~7d˰�ĕ/yF�����tuʵ�a�eHH��ƃk��)��b�f�4Ӛ��oy,]Ih�9��7�7���t)�p��a�L.���n��9Y���N���������Ri���@M��,���4�.b\ǲ�7P=���`�_��}f'oa�L>��'_��g���h�����Yb�!��T�����}�n�c'>�Է\�p�rA��\bxxc���ˬ��l�`@z.��.܍��G�e{sڤ�<I�ƻ}�b�S�u�t,8�s�ë?�nuV�|¸����|���sx�X:�Rݿɣg�NIA}�P�&�K�a����	�7E�ŝ����e��*�G�~�D)[ر��~<��4�ko�|1�A�ɥ_J���4�ͨ''�]&�F�'��?9���b��e��wWl�t'_T  f�i<��>�,]���oX���p�TA�D&O�{�t��I� U+��o��I�(�SMQ�'ׯ��r	m���G�PKRw0]Ok��Z2(���V:}�C��U����J�n_��G�i��*o�@N��xp}�mL!�X��'z������i�E���T-�J qAa͗t�/�/b~Z,�,`����_�;�Q �@��{�����Dx@�<T�G`��f��	O���K��]���LLL��yht
��z�֭9��������G���ҿ�u�M��_,8�M��^���i����/CɆ
�o��F���F�Nޠ��p���~0.7}��c��i�o�ې>��{=�qAW���^��x0���6���<�Kj����QM��q��Ҍ?X {+���{Y��z�sbr� �G^9E��۴ME�g�����>���K�w�fҍ/��AOt��M�F&�p$��u����L�����B��Ԗ�(2�����5w�.���ڴ�F�bW�O�Pe��}�F���F��&�<�L�1�!�X���_���U��ȓ�Tt�]��{[��L�FAL��� ^'��J�?���}��>Э��&T�uз�"~��US_�0��x���?N��]��o��o<d���>�ܺp�iS�#��nȗ8���dV	I����@g��\�����
\'eVJU�ە�;���D�а�����p_8���Hg������ƻr��U��5͓S̒� ��V�2s4U�����Pe
e�$"��]�#�.9���&a���:L�J!�/[��:<<%�$�׀ﱯˆ�^1͎��b��}�H��p5��Q�D�PIͥ�ݺ��U��_O�qz2�2��k�̏���|I��n_b��}p̓��.�����<.j.r�aX�Ic�>����K^��+��� ��b<�g�G��朗���0��s�ɭ���q\�q�IYQd���3YK��[����$�ڜ�{�I�!����i?b��s0���D�	@<m����Ĝ��R3����x��I)ehh9J�����U����e�H���&ш��q�{�%��ʠ��WՌT�!��*��,�O#ߙ��e4���|bGC-�!*糹���B��	��tV����k�b�.���
�������v߻'m�ԇ�&�K��3�x���g�n���`�]J�,
?���aMV���+��p,NP&���@�Gj4�7�(Ʒ������?��L�Ӷ	��ͯ��G������=R�ˮ8H�V=�����5\����:�
7�cXa'w�;�r�R���o;O����Y���V����߼6ݩ8؂W �7��)��v��y
.��e<h�p�ahISގ�2a�o�O�wDjjS�il��Q
 S����}D9h�C'�
���-}�L��\���2q�\)��I��*��`w@8�|F�po���gc��c���^\�>�����{��1q� ��M�zv����]�K���<�ŏpf��wM1$��%��f��u+��x��6����_�X���{ٔ%Ww�
y��A���P��j�dF�L��
�ֵ��hiM�~��CZ	c��n��N�k�V,��l	�'��3,��H�@�8�/��AǼ� �`�gb,� ���&��!�2k-� �0��*�8���]F�4q������(���ǘ=�ӊ���&��
����TY 2�B�KeQ���D�C�v���;9���ܒ��/��
s����.q���҄0��Ŗ��=+�=xD6N��=���)�&!T����O�|�l�v���!;͋��΅�EQmV�����U�ms0���Cs�e{I�:<KY�L�����;h�ؚyǜt��O<�������Bu�R-�_U'@"�q«j!�a�?\��+CFU�K�%G8@����A�h��8;��<�͜x1E�w�I�T$�Q����pz�%5��Jl����wU��wn�V��d���z&���zV�E��WI�iÂK; �ے�����w읢�@�
+e*��[uZ�п�T�R�4M�X�IY-����"G_#c�4�f�'�����Dg�I`�E���})�<�^g� �e�E���[���U�S��o`�v_�NÍ���YZЧ�Awס�W�b��p��0��E����;��U���(�"Qy�4ŝ(��7�z��%ha�gP+Ga���V[��;ĩ�%6{W����jy�jF{�B-���$TD���L���}��7�X��1�D����o��z�~-Z��1��A_�=li	�#t�J5)�Ph ����q�%r��7��*z��J��G�ߜ�0[\NOv�� ��0Qg0�\�<�v�)	����'Qא�E�QZ)P�^0&A�7u�h��'�Y]�Dʶ*�y��e����T��&�#qO�<����~��5�z����F7�7��9�����ʇ�>�@�a��B�1�Y������W*�M�a�n��( A�}PY�^�A���V` ��5a�7S���1�Fl=$�b����n�ǝ��ϝ����?�(��q�R�q�|N]c>I�{Ƒ�ԣ~�k���f��F�D�ڄ?hL�I6�{��Ѥ�5�,�]{4�H0��1��а�u<��C�D�qS�L;Pd�x�jT��,A�P23} <t]�J���6��x&ر~�XXnP�"�p��܍�p.<���MZ=l3��.��"	R	D�t���*�f*���g���Y��F��FO����F; j3$��]�Յ^��Gv#�B%0%�f`�#T.!(�¹�dS�切v����}��E!��,u����(�mp�F^��^�5�{������t��
��M�����qP>���:u�V�[�`�
���BE��U����L��Aنk'�Ӹgf9���6�jS1���s���ɪ7fp�0n`p��Գ���)j._��Ӧ���G�늊~�OT;%�:�BӇ�d���'s�	��?�וMA�x���';�|���U< �`
�%���g���"0��¹/���^���j�ó�k��ug���v/�9��أ�]���M1J"�5�����v���⏪��s�rn^PQ.�^^y��r���|ь�`	��(�^u���6wDZ��<\/bF��~��Ԡ �ᡛ.���WI�]�����g���Q�RË�Y���/	=�y&���'C�]�<[�TI�V� ƞ���~t�za����b�ꯦ"7�$���p$���DO��?�C��lR�]L�*��E��hL� i���e����}�w]�#���J�kw00��5,�f�6�5J�]7�D%���9�.-�fx�]�����Oa�JV[u��1I*a\+DٙPjUɆ��Q�*����O�:,�g- E�?�s�P1|�St1(�?�Ƭ5���^.b�s�_�;�gŷ�(�{/ -,K��f�xs����,	����vT�&[8��
��A���Z~V�M���v�Ō���\�1�Ӫr%�I9�}��tc����<�*p8�.���Vϔ[�ӵ���X�����Obӥ�v�υRU�]��̤{�:����C����L2:�r:�.:\���9֩������^�P����tV*=��s泂�#�/�#9�*Yl`�wuS��F���GNW'�ִ�"���Խ� ЙAH}�K�/ȅ��W3&f�7x"�J����I?�v�'��Yt�|'���O��
���A .٥�8?����LY �@�I��\�BU����B{B~�Hj{����P<�:P��>�nl�=2�i�b���2�#NU/����_�Ι*���7�\��Z��Cu���h�����ڕ
�\�٪�߳J�����%��M#�!��І��A�'��md�����Fu	�9�V3$�.�����"�}�F�a\������EPf��"lW-DL�b";�&d�2'�<�R�_�jM��/�k�S�-鉼�4�2LT��*�lˆ�it;����#�*�X�ײ��]���!\�vz�!"�Z�ȦI��Ɣ�Ƒ�"��
���}:I��7�(K8RA��N�Y�?@�x�a�Bvjp���-y�L�}U��gcJ�?��<���#�~�ZsA���Aru��	��S�C���#`^ou�kD�x��}A0�M�����O?�5�UL:����{HLŶ�����
&��0�������Ys�� w϶tpN�#��g�,�ŉ~n�����C�����)��������O|�i��94s�2_xک��Y���?]�a�z	e[��Aab��A�QMҵ'�k���ԑq/dY��`�WJ�_l95�K�^�{jz���DG4�2��l���(��j��-&b~�(F����r9�&"�&{��w�wA&/���׊�Laތh�v���!���3��RjM�D�����-i R�l$U[nkIB|��
"v���b;��0���t�;i���n(C�`��e�B�%���A�zZ2��-}d���R��H����![�}ʑ�g����&6���o�v1Fj�	Q���](����	�09����9�W����N�c�M�ϒ��y8g����2g$���Hq ��V��~�;�i���cљ?�-�l:;�d/�7Ga�a�L���_F�bJ@�[VB�Qr���,���7�ç����Bz/����1]lm��H���i��͂��E+:o|���ֻ��W���Z� �I�j
k�mcC�W�e�w�a��s�>���A����۾���0���b��	oS3����R�#WD��-˿o�ik"�"2K�K��=�޶R3k�=��Z��C�g6gY
��
[�@$ۦ�a����BU�k�$ê��\N6��,�g��L�=@�����[	�P-d���X�ϵ�����&��Ip�z��O�˥cŋ��C��}��xQ��c�`R�<�%C��)@�cB��*���@�4��Q]$���`v�6�-�vǊ�>�Ư�Vu
@���a����T�y��ٛ��Ѝ+�}��Axk�B�C�ܚ/O\zV:�i�99|��g���`�����(г�rHQigs��5m�z|Y_8BAa�F �S2�žT:��Q��-�g�1�K���������S; .,��t4`-26��7x�2���@X[���ߧZ�_U����Z���T[����C�3�V��:*�-�z��<���w��m��2����>�-������e,q�Z����޳��h�C�;''�l`G.�5#	D�)��"�q{���}c�pN��v�^����F�;A��\���w������ *�� J�3pb�BÒt�끪���&3SR�f0�J�Ԕ�팓Iʹ���ʉ�� P�v]�B(|bZo
�+iz3K�*k�Ӝ����әw{[��d�$L &+�\GP�S�����?�d�anz�"�~�5��X�QJLn��g���3͘7:oqə�������H�7���ix�����F�v���ɓf_��&W#��ڝ�@�?/�a豼�c�a32�=�[�ع��X���i$��qC	M|��C����#�˟��䏲՝`Mcx<g��R㊺1?�� �;���	�b�z}Fܡ���U3Z��1xq�b�i�G���8���n<_/�4�o�Ǿ;�Q.Ϝ8��gF�q>|Nu/m����6�94ը��	�l�\�8m&1g��|kHӾ��":`��DW FR�q��CoH�W��ݻ�<x��ai�Ex��b���~Fz
�� ���b�ey��Ϸd����e�,��&M���)@�sh�Pgn�6�-Tf�.��M�̉F"+l#�I���~X�3���X��P���m���8,NE���Z9�K�:o$�����N/=��%��(�c˗��[��X���QO2�0[Xqx�	����i/�~<���>����4�1Z澃`�*5�| tH�˿AzyC�L��[�S|�W��Wobu�������;!����5�T8��8��(�3]��e�����0k>�@X�l��k�2S?�ŻN6V'r�b�D��7�3���go�O��>h��Y�eJ�&�;�gvӸM|�* ��6 +���G�Mn�����p˂c�r�0!Ѡ3Hy�Y�\�]}�͙k(��-+Q�.� ��=ñ⫰�C*Q���öF&�0k��V}�:h�����M��'mEe]�"�N���w���E��$������9�bY��ɚr�?����s�s5���8�
S<�Fn���9��lB�rՎA�&u�L<;0a������ &�s�y�+�޶e��5֓B�8�ȋ>�)ցt��nr�\R��B5�zz��ɗ�u��3��	8�vj$�k� Q��W��2�Jm�U.��,{��u�N>$��h��5�b�<�^�b�>��)o& Q��{������[z/>2��1��V���:�,3.L�Î�1�Y]����Ҭ.��V����d�ӢG�E���S������_��t�P*�@G�sQq��  ��w�X�X۷8A�����>4m�a}�Dw����ދ��r�Г���V. 	�jK˘��M���Ϛ�'P*��m��T����4��:^XƾwN�o.��ϟ���Us�|���������f���
pu�=�J�D�N�y�g����W6��3����&�L�^�����οϨ�备�-Ze���|̣�Ϯ�Ś!R|�Aá����ې�c�'�}��9�ql��<̶�(�!r�;��6EZ�/��{�?j���Q.��	@���r�ʧ#��Y|����A�΍�w���Lv
@Y��s�S7E� ��H�� ��n]I:v� �h�Xt})�6�3Q`��
y�m�}�]M�b5�_��ۊ�*O�r$��k��9��'�O($����%�D�vm�c�k ـ�5[P��:d�I(&��ˀ|�rA%������z���g%}�D����Kh�����l��ec.zT��̥��L�E*zm��� ���l���!��"�{\G�������)@%}d��NC,�gb퐌h l�)?4Mn�`��K�xS���1��.}rKh�jՄ�ٽy��={䘪I�]1T��ʵ�D�����luF��/��NJ
c�(�� [Q��6_�ORg��*IT�'z6���Y�p =���)F~#�Lr�i��+����+��:���y��Z�d(�a7+��#ܤ�qٖ����z^��a=r�D�{}/��pg	�T$�\L�v;C`cӖ�e��7K�O�D�۴M��&�f��]��Y�2�>����LE���a`�}�c�<�7M��&�6����$h�χ��Z`�I� :/+@Bh�b�0;W�2ox�l'��������,k��]*p�g�h��PQtj�<���!4<���B���˷�*j���y#^[�����wίzO,Ar��D�Q�H���!�B��a�b�*u�Lלa�ߗ31}����T4�t����ӕG��S��G�F�(^@/W�ZoV�d	C�`�4��+�[]���r�"G]C����}o��F��[�0�먍X����� 8���᎘2�Pٶ�۪˴�?�<��;;�h�W���QV5��7��f��T5#�LU�v�1X^}S��T��z����
>�N�������
�
5���ƻc� �k�`p'`O[�W�B��qA��.�ɑ:mH�P��ҝI�{�uP#�A���˴��p��=I��-���D����/LX%ɻ�R�ev����((��1��R
��E>�IwN/'P�Qf3���</{p��Y����nSb(��=�� 9��"�)�C��<����a�Hd�i�@�@S=�P��j�V�����@wР	���x�_뼽R�\U������겅9g"Q8´��Ŭ�����1���{�*�T{gM���|�����݀x}�2�ޛ��d�A�+���2�%%ϳ��N5���^��kL�d?�bY���fbs\(ԝG���wxn��lΎݘ�KG�w�_9�ytS�cq���I{ܯ��h���e_	�>���nl��d�:�)���C;�$uԷm|�3��x��^<~�k�A~���h�ϭ�������u���#vE����b ��f��ZI,�ˌ�3�~�"��?9�<��Kf�IaiɒX���[7n�L��t@�`a�s�5g�Rk2��	i=��~�_[Ĕ�a�W�f��:��6>i8��Un;FY,%�Mg�np�9��H}������6����/�pp:��ǈ�����Vi�S��J���< o1�����k�L^�������p�N.Y�*3]��k�n����EV��;-�9)���7�{�3�W;���D�8�i
:�
�a�#�̖j�C^��?׾`��eT�uj���S������ܧ	�q��Rto�O���C��>	�>#�M��{�
b��N����H�(w&��f\ԋ3�ه���6��'�0�U�[���jV���G�8.B���Ĭ��֋�m2��R{���咓�%s��&:���G�`�P�|�����Rv��b���ID�Ӑ%���r/'P���mGp	'I��x�x�qν��"aÓ�4_��)�GR&�@TE9��-�{�%��S�ô���&f��j�N��%�����#�F_�:03���ի���?i����z�o����6��b�jB���)6)�i�6�빲0�Hľ����ѝy�Eu3���M�X��l��=�k1�U� 

jT��-|���4�9�.���3���d[�@��m:(�ϕ?��!��F\�-�%�b�YV {��.T�=v�����K��54�Pn��-��ժ�g�6�/��V藑D:K��{�~��dD.��֤���,Q��>���ή���'���^yB3s<����z�L�ā������� �w�[鶆������+q��ӴkbXU*U���[���?q�7�[�u�O����,���Eњ�19�á�< ���ة �ʻ��Vk��;8��]��=[��VR���r���e2s��)��z�~\C�Ⴈ'5�YАI���p�Av�/����h@ڽM��	s�^�܊�2@�-��ä�r1���p�&�X������GY'!�n��=<#�=u�ht�A�1#�-���0/8j3��˶�%�E�l���۞���N�b(��cU����Jm��s������{�͟@Z;�L4__Q$�
�6�t�����5��qk��ƾ&��n�	��I�k3,b#n�+�>�ܱ�7�CX��>�.x��(���7 ��K��k����;��q�GF�q"�$��`[fu{�dr��v�sՉ�����&��r�q�I��� ��Q���v�2�R_c�Z��JF�ѣ���a�9��7�(�֙ۉ2yY����-�VJ�(
��2F�r?�w	�$��5oI9�FFwI�T���CKx;����M��]K*��x�'���P�<�L���vj�@\��_�K:Y"��A�i�+�n�P��!s�gMX�Flu� ��f�	v���g�ӣX���
H{H,�d@�����	�P�J�;c�5U��Ւ���fw�E>��T�Y��7�-�G���^V�@���kdA�K%���0)r,[åv�9�;���ZM��J(l���(�����(4�Ehl�wQ���U#V���!��SmE��M�0W��{���3���<.�!J<�X2篼���%��ʰ�%��ß�XW��(e}@+����Ƣ�5�(���8�fxO��P�]{ּ�@����הG���8��ڐ�������c|Qٟ�(]R��_D9%t��ð�N��CvSXY�Ʌ5�T	�wG�xX<im�U�}�8,#���vdMG��{#hNAI;v���5q��yZܱ,+J7��G�e@(z�%G�P��@)]�k8+����k���dz;�׌�9e!d���Y����c�2���Ŋ�� �4�J+�,��X��z�f�ӢR@�0O�*���|?[�#6���4Xj��r;0
�:"�-��h;K<":�	�+��Cr[qq�m��T�MM���K�:�ڱ���RY���t��` w��פ�Ԯ�
��l�ɮ����*MlV���k�`�$���t[��3:��ˁY�Y��T�u��[���nl|�9�١=�W�NU�|3�뫷6��i�߬�����P��Q� :��փS��Q�����g.��x�ǳ���������ז�s�Q$�q��6I��lB��y��7�}~�k�gmm\�/{�q]i����� I�Z�s�RY	���G�\��G�ُYy�V,ߺv12�9�=���)c����drx�C������
����L�B�3-)+�t_ʅ�_�-�7��J@��S�����ο�a��aF?��!˕� �9Z��!������Mlһ�㳏����)��4K��	oVND��B߭�3��L��2o�]���G>�^��d�Ӱ�VU�MF�����=3�˚���-�x;�6	���n�ӓGU�����|��b�ꈵ��A扄9b�����>C�3ρUD�d@+r���o��B�G����s7�C�e�M��d��׫�.V�)1�����\�~���w
��:���Rb��B-��U����D���v>�r�xMB�y���1�z�,�^��,���<�G�x�u�m�Ϋ`=�2=ti��[e w�dt"<�i�� �&����_��㐐��u�%�N?���>�G&�E�qHy����C��N���1����u�N�Ԉ���Y���ʳ:�����t�j�ps`/A�/���O�ta�y�H����bPه�{6���k��~� L�;,	�wpv�>�pc��cQ����UJW��'+�a�K�-����?�SMy���V5�j@�<-��BWo;��"�to�oA�ݓ��a,�[�P�$�{�eb�\�Zڕ����p����oMaQ�s�nt�Z2g+]2 �|��*D8-������uH,���5�˷�޸�T�0%O�E; �Oi�5p��.��P�E�ػ㥢H]�x����Fρ+����s?�ލ���g��;�k��	5�r�S��-�`���8}<o/���sd�����"�P�T<�� �pz̀6�q��(�p��9�}\�2��\�}���a�:5��\՜Z�p(��K�e�1s�����"^���*ɟP����E�3PJSK���~yJ�t��C@�6HB�j�o(CI�N�A���Lki/�Ļ�3�6z����vX��k��²Ǣw5���Ronu�=kDai�F��ic{wc/s.x=�C1h���hOe�[��J��	���W�22��,����ȗ�y[����5Me�!q�z���L kLP	N���������ٿ�-j��"C5I�;\ B��[�bR����Ԅc�S�;*���Ɣ�Y#���ѣ�Th-�g��RC�� f��vT�$���x���݌E��$�\)�3΢�'��磄b��J�'��,E�@*Y�I����LF��ɶ�u��r!�j]m�����*_r��ƞ^@��� ��8P'
�Z^�0_q۽��K���ERP�)o�n���������J�V0$���g"}~M����0�y_�
�^�}�F�Z[%W<̌86u�MM�V�4���!<z�zH�#?o8��J灻�C	�rw�Y�w���f��%C'�l �B�d���֎v�Y�(����m��_�08���ʼt�����#���p�\m[E^�r�%*j� �N��"����k��y"�o�h[B�����.��P��T�XX����|�>���~��m����H~���Ĺ�L����<�3�o�w�q�̠�Nl`��Y��ȶ|��8%�9X�K:Jd��'�e�Rqř4ȋt��%�jΝ�����=|/(�����1@�,S��6jD/��wv�oT_��PL<�h�z�uu�2�-���}��Z漑R5h�����!]�G��@�J��؀�?�,��L��!1�4]
�0���X9��z f&Y%���1�לr�N�y���T��VtW����'��M6����M�ك�Q7`�(��tf��_�<�˰�F���p���9a �ޏ6b_1���8s�3��j��m���t?�ɉVO�KA��0f~���x�"��C��nQU���I�'�zC��nH!h��åM��������bDe�%�G�n��a3�AX�e�AI��|oMe�ں���\�����������=H<\�f���i�����Pj��>%@��R������>y�T��Y�͉�ܔ�spD������ˁp��ə+�3�Z��@f�z焫[��0o����d�
,�"{���ˊ��ؚz������Q�����f��%�M�d,ҽ;&�e>�	"{?#��j�0]��c.9P�3��<����kR���b��Z��x^�=�&M	z/�$��d�"J���B, J�s��M.J¯���A�g܃���Y9Hl�N����&I��oγ����u�md�\�9�.J-��&�+>�Ǐ�W�i�7��B��o���lu-�U:j2��(L���൓���SJVt�)��j uZr�o�ಅ�h	=Z[���r��o� ����H�s{���G�8���y��h��/,�"�r����b�UYb3�Vcݱ�ZX�X�V���w��kj����9�����R�i���[���݁_?�&�Y���v��n����k1�qrթ��Od�����"�G)	��s���y
��s��&$}l�Y���?De��*�6�������3�V.|PJ�W��z^�-��`i=Ĺ����fG��!�����1�*Б����=��&%o���y 10R�U�&���q�ec`��4�V#�A�Zҙv��Vw�Y���#��y���C��k�9���A4�,���@�ƪ6ޯ9 S�M�H��sp{����g�>EY!�c���0kd/^?W���r�����>$�D^\�}PC���_H(R��JiX�֮f&��9�j��_uS<�Ĉ<IaYE�!2�qP5��.[D��*;Jd���fV��c�,�ۏQ KK�i牎d��_�i�4O&R+_T�?��� "9��{�-B_�{7�P �
u�	`�C�����^��a�*Uђ��K��R}J�ф�s�K����~(;�Q�LEC}�Gg��+�C�%Cg����o~�'Od��hH߹^Ǖ+9e��K�8�(��R�7�U�[.������FηN�[ �I0�[���8�����	7�ѫqJ�O3Gq�ڡ��y����u��@gg���z��Ŷƃ .}�hĞN<���-V�-w��$���#X��I���&�Ñ�c����YԖ�T&I�_��pu�_rꭀ`���j^�.�ks� �o����7��[�ԓ��G�Q�)y[�����Y�٫�ry��(W+;,w����*N���c�Y��~Ե߯��Q����]���m���%\�T���<��ɒb�Z�P7�HW�a�ʂ@����ڍ0����>�-~��	�zm9�W�U��k�ѯ�e�;����U �?-�Y���cs���1�=��ۅ[�b/j�u����󷭩j�Y�ꟸM��� ���?T��%���>G���Ɇ�^�����/:�%��]��0"�%�2�,F�*� ?���,�@����y��|�;������U�ީ��Zp�%Ѻ79�ڨ4^��q�: 	R�?��^���=��P�FV
~�kA˃r���M�'�p�;�$Q�Ȭ�YT<�W�=ؔEuԢ7tEȓ��D.��Y��h�Zs�X��?�X�?���/�)����.�r���߷��b��d[��/��ǖ�A�|$�6:��v����s�/hj6a�� ����\��	�5�?�/5Qt�	*lN�h��)��Ei��Rr�ƙPɏu��l~�o8�0�C҄8	�M��p�AHp�����bU9�����Kv� K~=��n�D�g��� ���Q�a����l�][���T��1��i�Nw8趱g�g�H�����݋�*�����?�F?��z(<�4��Xz��Z-�s���47ysa�0A>�z����zI��PL��bN������1�h�1`���ѩ`�����Ub�/�z\%R�WE�׶�uǮ{�15Tc��@��+ ��w�������&X*S@䙕3��z��l����E�W9�F�X4�Y �}��r��k�t�$2��?�=�8�r�=UQ�6{Hfa�(���=���{j*XG��=�@��×�)�`�W�6 �{�H�f��ٻ!I��o���ďC{/�3��X)��C�9������������:
�"��1i*�,�lX �ـ�{��t, ��T2f���V/Ua6��9����|7F�:xL�\U-�,�0Q�������'�ԮF}�P6���4{w��!�Q�s̲�k�N�E�=���jj5Y�_����(�e�!���lx:8.i�/ufĮ���ar���C��{P iG����"L�B���Z.D�}�]�ty��9���b*�J;,s}����\�����
��o��_�u$;��>�4L��=����=�P,�����Rǝ/$��N�4��T�zA���ƎZ��v��X��y=�������R����r5�������.����*&Ϫi�ݽ���9�H�������)�)�˲�έ��,��Vo0�u�#�J/�0u5�q�㒷iI��f�P��L�����P���gl��?F>������M~`�e�Hc��;��q?%L҅��[��Ve�ҧ���G��y��信�|s��y	�����Q���ԱviцE�t��4���1���#�[~�%�!�ϑ?� �S�8z.۶g����q5�w�j1Ml2!��K�D���J����u�9�*B����C�f