    Mac OS X            	   2   �     +                                      ATTR      +   �   o                  �   S  com.dropbox.attributes          com.dropbox.attrs    x��VJ)�/Hʯ�O��I�L���ON�Q�R�V�ML����%����RK���|߈��L�4���0�2Ϫ*3o�t[[���Z ͜�

�!�WJ>�     wD��ڞ